`ifndef INITIAL_DOODLE_LEFT

// Module definition:
// logic [79:0][79:0][2:0][3:0] doodle_left_rgb;
// logic [79:0][79:0] doodle_left_alpha;

`define INITIAL_DOODLE_LEFT \
always_comb begin \
	doodle_left_rgb[0][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[0][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[1][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[2][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[3][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[4][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[5][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[6][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[7][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[8][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[9][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[10][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[11][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[12][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[13][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[14][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[15][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[16][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[17][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[18][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[19][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[20][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[20][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[21][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[21][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[22][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[22][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[23][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[23][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[24][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[24][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[25][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[25][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[26][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[26][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[27][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[27][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[28][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[28][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[29][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[29][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[30][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[30][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[31][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[31][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[32][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[32][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[33][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[33][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[34][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[34][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[35][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[35][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[36][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[36][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[37][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[37][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][8] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][9] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][10] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][11] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][16] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][17] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][18] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][19] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][20] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][21] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][22] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][23] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][24] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][25] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][26] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[38][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[38][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][8] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][9] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][10] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][11] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][16] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][17] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][18] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][19] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][20] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][21] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][22] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][23] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][24] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][25] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][26] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[39][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[39][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][8] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][9] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][10] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][11] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][16] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][17] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][18] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][19] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][20] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][21] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][22] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][23] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][24] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][25] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][26] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[40][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[40][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][8] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][9] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][10] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][11] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][16] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][17] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][18] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][19] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][20] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][21] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][22] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][23] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][24] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][25] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][26] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[41][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[41][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[42][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[42][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[43][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[43][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[44][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[44][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[45][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[45][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[46][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[46][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[47][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[47][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[48][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[48][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[49][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[49][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[50][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[50][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[51][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[51][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[52][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[53][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[54][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[55][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[56][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[56][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[57][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[57][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[58][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[58][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[59][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[59][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[60][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[60][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[61][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[61][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[62][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[62][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][27] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][28] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][29] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][30] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][31] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][32] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][33] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][34] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][35] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][36] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][37] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][38] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][39] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][40] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][41] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][42] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][43] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][44] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][45] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][46] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][47] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][48] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][49] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][50] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][51] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][52] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][53] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][54] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][55] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][56] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][57] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][58] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][59] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][60] = {4'b0, 4'b1111, 4'b0}; \
	doodle_left_rgb[63][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[63][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[64][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[65][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[66][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[67][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[68][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[69][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[70][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[71][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[72][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[73][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[74][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[75][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[76][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[77][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[78][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][0] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][1] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][2] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][3] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][4] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][5] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][6] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][7] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][8] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][9] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][10] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][11] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][12] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][13] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][14] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][15] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][16] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][17] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][18] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][19] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][20] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][21] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][22] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][23] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][24] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][25] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][26] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][27] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][28] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][29] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][30] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][31] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][32] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][33] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][34] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][35] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][36] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][37] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][38] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][39] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][40] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][41] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][42] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][43] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][44] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][45] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][46] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][47] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][48] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][49] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][50] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][51] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][52] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][53] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][54] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][55] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][56] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][57] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][58] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][59] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][60] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][61] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][62] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][63] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][64] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][65] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][66] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][67] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][68] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][69] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][70] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][71] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][72] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][73] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][74] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][75] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][76] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][77] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][78] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_rgb[79][79] = {4'b0, 4'b0, 4'b0}; \
	doodle_left_alpha[0][0] = 1'b1; \
	doodle_left_alpha[0][1] = 1'b1; \
	doodle_left_alpha[0][2] = 1'b1; \
	doodle_left_alpha[0][3] = 1'b1; \
	doodle_left_alpha[0][4] = 1'b1; \
	doodle_left_alpha[0][5] = 1'b1; \
	doodle_left_alpha[0][6] = 1'b1; \
	doodle_left_alpha[0][7] = 1'b1; \
	doodle_left_alpha[0][8] = 1'b1; \
	doodle_left_alpha[0][9] = 1'b1; \
	doodle_left_alpha[0][10] = 1'b1; \
	doodle_left_alpha[0][11] = 1'b1; \
	doodle_left_alpha[0][12] = 1'b1; \
	doodle_left_alpha[0][13] = 1'b1; \
	doodle_left_alpha[0][14] = 1'b1; \
	doodle_left_alpha[0][15] = 1'b1; \
	doodle_left_alpha[0][16] = 1'b1; \
	doodle_left_alpha[0][17] = 1'b1; \
	doodle_left_alpha[0][18] = 1'b1; \
	doodle_left_alpha[0][19] = 1'b1; \
	doodle_left_alpha[0][20] = 1'b1; \
	doodle_left_alpha[0][21] = 1'b1; \
	doodle_left_alpha[0][22] = 1'b1; \
	doodle_left_alpha[0][23] = 1'b1; \
	doodle_left_alpha[0][24] = 1'b1; \
	doodle_left_alpha[0][25] = 1'b1; \
	doodle_left_alpha[0][26] = 1'b1; \
	doodle_left_alpha[0][27] = 1'b1; \
	doodle_left_alpha[0][28] = 1'b1; \
	doodle_left_alpha[0][29] = 1'b1; \
	doodle_left_alpha[0][30] = 1'b1; \
	doodle_left_alpha[0][31] = 1'b1; \
	doodle_left_alpha[0][32] = 1'b1; \
	doodle_left_alpha[0][33] = 1'b1; \
	doodle_left_alpha[0][34] = 1'b1; \
	doodle_left_alpha[0][35] = 1'b1; \
	doodle_left_alpha[0][36] = 1'b1; \
	doodle_left_alpha[0][37] = 1'b1; \
	doodle_left_alpha[0][38] = 1'b1; \
	doodle_left_alpha[0][39] = 1'b1; \
	doodle_left_alpha[0][40] = 1'b1; \
	doodle_left_alpha[0][41] = 1'b1; \
	doodle_left_alpha[0][42] = 1'b1; \
	doodle_left_alpha[0][43] = 1'b1; \
	doodle_left_alpha[0][44] = 1'b1; \
	doodle_left_alpha[0][45] = 1'b1; \
	doodle_left_alpha[0][46] = 1'b1; \
	doodle_left_alpha[0][47] = 1'b1; \
	doodle_left_alpha[0][48] = 1'b1; \
	doodle_left_alpha[0][49] = 1'b1; \
	doodle_left_alpha[0][50] = 1'b1; \
	doodle_left_alpha[0][51] = 1'b1; \
	doodle_left_alpha[0][52] = 1'b1; \
	doodle_left_alpha[0][53] = 1'b1; \
	doodle_left_alpha[0][54] = 1'b1; \
	doodle_left_alpha[0][55] = 1'b1; \
	doodle_left_alpha[0][56] = 1'b1; \
	doodle_left_alpha[0][57] = 1'b1; \
	doodle_left_alpha[0][58] = 1'b1; \
	doodle_left_alpha[0][59] = 1'b1; \
	doodle_left_alpha[0][60] = 1'b1; \
	doodle_left_alpha[0][61] = 1'b1; \
	doodle_left_alpha[0][62] = 1'b1; \
	doodle_left_alpha[0][63] = 1'b1; \
	doodle_left_alpha[0][64] = 1'b1; \
	doodle_left_alpha[0][65] = 1'b1; \
	doodle_left_alpha[0][66] = 1'b1; \
	doodle_left_alpha[0][67] = 1'b1; \
	doodle_left_alpha[0][68] = 1'b1; \
	doodle_left_alpha[0][69] = 1'b1; \
	doodle_left_alpha[0][70] = 1'b1; \
	doodle_left_alpha[0][71] = 1'b1; \
	doodle_left_alpha[0][72] = 1'b1; \
	doodle_left_alpha[0][73] = 1'b1; \
	doodle_left_alpha[0][74] = 1'b1; \
	doodle_left_alpha[0][75] = 1'b1; \
	doodle_left_alpha[0][76] = 1'b1; \
	doodle_left_alpha[0][77] = 1'b1; \
	doodle_left_alpha[0][78] = 1'b1; \
	doodle_left_alpha[0][79] = 1'b1; \
	doodle_left_alpha[1][0] = 1'b1; \
	doodle_left_alpha[1][1] = 1'b1; \
	doodle_left_alpha[1][2] = 1'b1; \
	doodle_left_alpha[1][3] = 1'b1; \
	doodle_left_alpha[1][4] = 1'b1; \
	doodle_left_alpha[1][5] = 1'b1; \
	doodle_left_alpha[1][6] = 1'b1; \
	doodle_left_alpha[1][7] = 1'b1; \
	doodle_left_alpha[1][8] = 1'b1; \
	doodle_left_alpha[1][9] = 1'b1; \
	doodle_left_alpha[1][10] = 1'b1; \
	doodle_left_alpha[1][11] = 1'b1; \
	doodle_left_alpha[1][12] = 1'b1; \
	doodle_left_alpha[1][13] = 1'b1; \
	doodle_left_alpha[1][14] = 1'b1; \
	doodle_left_alpha[1][15] = 1'b1; \
	doodle_left_alpha[1][16] = 1'b1; \
	doodle_left_alpha[1][17] = 1'b1; \
	doodle_left_alpha[1][18] = 1'b1; \
	doodle_left_alpha[1][19] = 1'b1; \
	doodle_left_alpha[1][20] = 1'b1; \
	doodle_left_alpha[1][21] = 1'b1; \
	doodle_left_alpha[1][22] = 1'b1; \
	doodle_left_alpha[1][23] = 1'b1; \
	doodle_left_alpha[1][24] = 1'b1; \
	doodle_left_alpha[1][25] = 1'b1; \
	doodle_left_alpha[1][26] = 1'b1; \
	doodle_left_alpha[1][27] = 1'b1; \
	doodle_left_alpha[1][28] = 1'b1; \
	doodle_left_alpha[1][29] = 1'b1; \
	doodle_left_alpha[1][30] = 1'b1; \
	doodle_left_alpha[1][31] = 1'b1; \
	doodle_left_alpha[1][32] = 1'b1; \
	doodle_left_alpha[1][33] = 1'b1; \
	doodle_left_alpha[1][34] = 1'b1; \
	doodle_left_alpha[1][35] = 1'b1; \
	doodle_left_alpha[1][36] = 1'b1; \
	doodle_left_alpha[1][37] = 1'b1; \
	doodle_left_alpha[1][38] = 1'b1; \
	doodle_left_alpha[1][39] = 1'b1; \
	doodle_left_alpha[1][40] = 1'b1; \
	doodle_left_alpha[1][41] = 1'b1; \
	doodle_left_alpha[1][42] = 1'b1; \
	doodle_left_alpha[1][43] = 1'b1; \
	doodle_left_alpha[1][44] = 1'b1; \
	doodle_left_alpha[1][45] = 1'b1; \
	doodle_left_alpha[1][46] = 1'b1; \
	doodle_left_alpha[1][47] = 1'b1; \
	doodle_left_alpha[1][48] = 1'b1; \
	doodle_left_alpha[1][49] = 1'b1; \
	doodle_left_alpha[1][50] = 1'b1; \
	doodle_left_alpha[1][51] = 1'b1; \
	doodle_left_alpha[1][52] = 1'b1; \
	doodle_left_alpha[1][53] = 1'b1; \
	doodle_left_alpha[1][54] = 1'b1; \
	doodle_left_alpha[1][55] = 1'b1; \
	doodle_left_alpha[1][56] = 1'b1; \
	doodle_left_alpha[1][57] = 1'b1; \
	doodle_left_alpha[1][58] = 1'b1; \
	doodle_left_alpha[1][59] = 1'b1; \
	doodle_left_alpha[1][60] = 1'b1; \
	doodle_left_alpha[1][61] = 1'b1; \
	doodle_left_alpha[1][62] = 1'b1; \
	doodle_left_alpha[1][63] = 1'b1; \
	doodle_left_alpha[1][64] = 1'b1; \
	doodle_left_alpha[1][65] = 1'b1; \
	doodle_left_alpha[1][66] = 1'b1; \
	doodle_left_alpha[1][67] = 1'b1; \
	doodle_left_alpha[1][68] = 1'b1; \
	doodle_left_alpha[1][69] = 1'b1; \
	doodle_left_alpha[1][70] = 1'b1; \
	doodle_left_alpha[1][71] = 1'b1; \
	doodle_left_alpha[1][72] = 1'b1; \
	doodle_left_alpha[1][73] = 1'b1; \
	doodle_left_alpha[1][74] = 1'b1; \
	doodle_left_alpha[1][75] = 1'b1; \
	doodle_left_alpha[1][76] = 1'b1; \
	doodle_left_alpha[1][77] = 1'b1; \
	doodle_left_alpha[1][78] = 1'b1; \
	doodle_left_alpha[1][79] = 1'b1; \
	doodle_left_alpha[2][0] = 1'b1; \
	doodle_left_alpha[2][1] = 1'b1; \
	doodle_left_alpha[2][2] = 1'b1; \
	doodle_left_alpha[2][3] = 1'b1; \
	doodle_left_alpha[2][4] = 1'b1; \
	doodle_left_alpha[2][5] = 1'b1; \
	doodle_left_alpha[2][6] = 1'b1; \
	doodle_left_alpha[2][7] = 1'b1; \
	doodle_left_alpha[2][8] = 1'b1; \
	doodle_left_alpha[2][9] = 1'b1; \
	doodle_left_alpha[2][10] = 1'b1; \
	doodle_left_alpha[2][11] = 1'b1; \
	doodle_left_alpha[2][12] = 1'b1; \
	doodle_left_alpha[2][13] = 1'b1; \
	doodle_left_alpha[2][14] = 1'b1; \
	doodle_left_alpha[2][15] = 1'b1; \
	doodle_left_alpha[2][16] = 1'b1; \
	doodle_left_alpha[2][17] = 1'b1; \
	doodle_left_alpha[2][18] = 1'b1; \
	doodle_left_alpha[2][19] = 1'b1; \
	doodle_left_alpha[2][20] = 1'b1; \
	doodle_left_alpha[2][21] = 1'b1; \
	doodle_left_alpha[2][22] = 1'b1; \
	doodle_left_alpha[2][23] = 1'b1; \
	doodle_left_alpha[2][24] = 1'b1; \
	doodle_left_alpha[2][25] = 1'b1; \
	doodle_left_alpha[2][26] = 1'b1; \
	doodle_left_alpha[2][27] = 1'b1; \
	doodle_left_alpha[2][28] = 1'b1; \
	doodle_left_alpha[2][29] = 1'b1; \
	doodle_left_alpha[2][30] = 1'b1; \
	doodle_left_alpha[2][31] = 1'b1; \
	doodle_left_alpha[2][32] = 1'b1; \
	doodle_left_alpha[2][33] = 1'b1; \
	doodle_left_alpha[2][34] = 1'b1; \
	doodle_left_alpha[2][35] = 1'b1; \
	doodle_left_alpha[2][36] = 1'b1; \
	doodle_left_alpha[2][37] = 1'b1; \
	doodle_left_alpha[2][38] = 1'b1; \
	doodle_left_alpha[2][39] = 1'b1; \
	doodle_left_alpha[2][40] = 1'b1; \
	doodle_left_alpha[2][41] = 1'b1; \
	doodle_left_alpha[2][42] = 1'b1; \
	doodle_left_alpha[2][43] = 1'b1; \
	doodle_left_alpha[2][44] = 1'b1; \
	doodle_left_alpha[2][45] = 1'b1; \
	doodle_left_alpha[2][46] = 1'b1; \
	doodle_left_alpha[2][47] = 1'b1; \
	doodle_left_alpha[2][48] = 1'b1; \
	doodle_left_alpha[2][49] = 1'b1; \
	doodle_left_alpha[2][50] = 1'b1; \
	doodle_left_alpha[2][51] = 1'b1; \
	doodle_left_alpha[2][52] = 1'b1; \
	doodle_left_alpha[2][53] = 1'b1; \
	doodle_left_alpha[2][54] = 1'b1; \
	doodle_left_alpha[2][55] = 1'b1; \
	doodle_left_alpha[2][56] = 1'b1; \
	doodle_left_alpha[2][57] = 1'b1; \
	doodle_left_alpha[2][58] = 1'b1; \
	doodle_left_alpha[2][59] = 1'b1; \
	doodle_left_alpha[2][60] = 1'b1; \
	doodle_left_alpha[2][61] = 1'b1; \
	doodle_left_alpha[2][62] = 1'b1; \
	doodle_left_alpha[2][63] = 1'b1; \
	doodle_left_alpha[2][64] = 1'b1; \
	doodle_left_alpha[2][65] = 1'b1; \
	doodle_left_alpha[2][66] = 1'b1; \
	doodle_left_alpha[2][67] = 1'b1; \
	doodle_left_alpha[2][68] = 1'b1; \
	doodle_left_alpha[2][69] = 1'b1; \
	doodle_left_alpha[2][70] = 1'b1; \
	doodle_left_alpha[2][71] = 1'b1; \
	doodle_left_alpha[2][72] = 1'b1; \
	doodle_left_alpha[2][73] = 1'b1; \
	doodle_left_alpha[2][74] = 1'b1; \
	doodle_left_alpha[2][75] = 1'b1; \
	doodle_left_alpha[2][76] = 1'b1; \
	doodle_left_alpha[2][77] = 1'b1; \
	doodle_left_alpha[2][78] = 1'b1; \
	doodle_left_alpha[2][79] = 1'b1; \
	doodle_left_alpha[3][0] = 1'b1; \
	doodle_left_alpha[3][1] = 1'b1; \
	doodle_left_alpha[3][2] = 1'b1; \
	doodle_left_alpha[3][3] = 1'b1; \
	doodle_left_alpha[3][4] = 1'b1; \
	doodle_left_alpha[3][5] = 1'b1; \
	doodle_left_alpha[3][6] = 1'b1; \
	doodle_left_alpha[3][7] = 1'b1; \
	doodle_left_alpha[3][8] = 1'b1; \
	doodle_left_alpha[3][9] = 1'b1; \
	doodle_left_alpha[3][10] = 1'b1; \
	doodle_left_alpha[3][11] = 1'b1; \
	doodle_left_alpha[3][12] = 1'b1; \
	doodle_left_alpha[3][13] = 1'b1; \
	doodle_left_alpha[3][14] = 1'b1; \
	doodle_left_alpha[3][15] = 1'b1; \
	doodle_left_alpha[3][16] = 1'b1; \
	doodle_left_alpha[3][17] = 1'b1; \
	doodle_left_alpha[3][18] = 1'b1; \
	doodle_left_alpha[3][19] = 1'b1; \
	doodle_left_alpha[3][20] = 1'b1; \
	doodle_left_alpha[3][21] = 1'b1; \
	doodle_left_alpha[3][22] = 1'b1; \
	doodle_left_alpha[3][23] = 1'b1; \
	doodle_left_alpha[3][24] = 1'b1; \
	doodle_left_alpha[3][25] = 1'b1; \
	doodle_left_alpha[3][26] = 1'b1; \
	doodle_left_alpha[3][27] = 1'b1; \
	doodle_left_alpha[3][28] = 1'b1; \
	doodle_left_alpha[3][29] = 1'b1; \
	doodle_left_alpha[3][30] = 1'b1; \
	doodle_left_alpha[3][31] = 1'b1; \
	doodle_left_alpha[3][32] = 1'b1; \
	doodle_left_alpha[3][33] = 1'b1; \
	doodle_left_alpha[3][34] = 1'b1; \
	doodle_left_alpha[3][35] = 1'b1; \
	doodle_left_alpha[3][36] = 1'b1; \
	doodle_left_alpha[3][37] = 1'b1; \
	doodle_left_alpha[3][38] = 1'b1; \
	doodle_left_alpha[3][39] = 1'b1; \
	doodle_left_alpha[3][40] = 1'b1; \
	doodle_left_alpha[3][41] = 1'b1; \
	doodle_left_alpha[3][42] = 1'b1; \
	doodle_left_alpha[3][43] = 1'b1; \
	doodle_left_alpha[3][44] = 1'b1; \
	doodle_left_alpha[3][45] = 1'b1; \
	doodle_left_alpha[3][46] = 1'b1; \
	doodle_left_alpha[3][47] = 1'b1; \
	doodle_left_alpha[3][48] = 1'b1; \
	doodle_left_alpha[3][49] = 1'b1; \
	doodle_left_alpha[3][50] = 1'b1; \
	doodle_left_alpha[3][51] = 1'b1; \
	doodle_left_alpha[3][52] = 1'b1; \
	doodle_left_alpha[3][53] = 1'b1; \
	doodle_left_alpha[3][54] = 1'b1; \
	doodle_left_alpha[3][55] = 1'b1; \
	doodle_left_alpha[3][56] = 1'b1; \
	doodle_left_alpha[3][57] = 1'b1; \
	doodle_left_alpha[3][58] = 1'b1; \
	doodle_left_alpha[3][59] = 1'b1; \
	doodle_left_alpha[3][60] = 1'b1; \
	doodle_left_alpha[3][61] = 1'b1; \
	doodle_left_alpha[3][62] = 1'b1; \
	doodle_left_alpha[3][63] = 1'b1; \
	doodle_left_alpha[3][64] = 1'b1; \
	doodle_left_alpha[3][65] = 1'b1; \
	doodle_left_alpha[3][66] = 1'b1; \
	doodle_left_alpha[3][67] = 1'b1; \
	doodle_left_alpha[3][68] = 1'b1; \
	doodle_left_alpha[3][69] = 1'b1; \
	doodle_left_alpha[3][70] = 1'b1; \
	doodle_left_alpha[3][71] = 1'b1; \
	doodle_left_alpha[3][72] = 1'b1; \
	doodle_left_alpha[3][73] = 1'b1; \
	doodle_left_alpha[3][74] = 1'b1; \
	doodle_left_alpha[3][75] = 1'b1; \
	doodle_left_alpha[3][76] = 1'b1; \
	doodle_left_alpha[3][77] = 1'b1; \
	doodle_left_alpha[3][78] = 1'b1; \
	doodle_left_alpha[3][79] = 1'b1; \
	doodle_left_alpha[4][0] = 1'b1; \
	doodle_left_alpha[4][1] = 1'b1; \
	doodle_left_alpha[4][2] = 1'b1; \
	doodle_left_alpha[4][3] = 1'b1; \
	doodle_left_alpha[4][4] = 1'b1; \
	doodle_left_alpha[4][5] = 1'b1; \
	doodle_left_alpha[4][6] = 1'b1; \
	doodle_left_alpha[4][7] = 1'b1; \
	doodle_left_alpha[4][8] = 1'b1; \
	doodle_left_alpha[4][9] = 1'b1; \
	doodle_left_alpha[4][10] = 1'b1; \
	doodle_left_alpha[4][11] = 1'b1; \
	doodle_left_alpha[4][12] = 1'b1; \
	doodle_left_alpha[4][13] = 1'b1; \
	doodle_left_alpha[4][14] = 1'b1; \
	doodle_left_alpha[4][15] = 1'b1; \
	doodle_left_alpha[4][16] = 1'b1; \
	doodle_left_alpha[4][17] = 1'b1; \
	doodle_left_alpha[4][18] = 1'b1; \
	doodle_left_alpha[4][19] = 1'b1; \
	doodle_left_alpha[4][20] = 1'b1; \
	doodle_left_alpha[4][21] = 1'b1; \
	doodle_left_alpha[4][22] = 1'b1; \
	doodle_left_alpha[4][23] = 1'b1; \
	doodle_left_alpha[4][24] = 1'b1; \
	doodle_left_alpha[4][25] = 1'b1; \
	doodle_left_alpha[4][26] = 1'b1; \
	doodle_left_alpha[4][27] = 1'b1; \
	doodle_left_alpha[4][28] = 1'b1; \
	doodle_left_alpha[4][29] = 1'b1; \
	doodle_left_alpha[4][30] = 1'b1; \
	doodle_left_alpha[4][31] = 1'b1; \
	doodle_left_alpha[4][32] = 1'b1; \
	doodle_left_alpha[4][33] = 1'b1; \
	doodle_left_alpha[4][34] = 1'b1; \
	doodle_left_alpha[4][35] = 1'b1; \
	doodle_left_alpha[4][36] = 1'b1; \
	doodle_left_alpha[4][37] = 1'b1; \
	doodle_left_alpha[4][38] = 1'b1; \
	doodle_left_alpha[4][39] = 1'b1; \
	doodle_left_alpha[4][40] = 1'b1; \
	doodle_left_alpha[4][41] = 1'b1; \
	doodle_left_alpha[4][42] = 1'b1; \
	doodle_left_alpha[4][43] = 1'b1; \
	doodle_left_alpha[4][44] = 1'b1; \
	doodle_left_alpha[4][45] = 1'b1; \
	doodle_left_alpha[4][46] = 1'b1; \
	doodle_left_alpha[4][47] = 1'b1; \
	doodle_left_alpha[4][48] = 1'b1; \
	doodle_left_alpha[4][49] = 1'b1; \
	doodle_left_alpha[4][50] = 1'b1; \
	doodle_left_alpha[4][51] = 1'b1; \
	doodle_left_alpha[4][52] = 1'b1; \
	doodle_left_alpha[4][53] = 1'b1; \
	doodle_left_alpha[4][54] = 1'b1; \
	doodle_left_alpha[4][55] = 1'b1; \
	doodle_left_alpha[4][56] = 1'b1; \
	doodle_left_alpha[4][57] = 1'b1; \
	doodle_left_alpha[4][58] = 1'b1; \
	doodle_left_alpha[4][59] = 1'b1; \
	doodle_left_alpha[4][60] = 1'b1; \
	doodle_left_alpha[4][61] = 1'b1; \
	doodle_left_alpha[4][62] = 1'b1; \
	doodle_left_alpha[4][63] = 1'b1; \
	doodle_left_alpha[4][64] = 1'b1; \
	doodle_left_alpha[4][65] = 1'b1; \
	doodle_left_alpha[4][66] = 1'b1; \
	doodle_left_alpha[4][67] = 1'b1; \
	doodle_left_alpha[4][68] = 1'b1; \
	doodle_left_alpha[4][69] = 1'b1; \
	doodle_left_alpha[4][70] = 1'b1; \
	doodle_left_alpha[4][71] = 1'b1; \
	doodle_left_alpha[4][72] = 1'b1; \
	doodle_left_alpha[4][73] = 1'b1; \
	doodle_left_alpha[4][74] = 1'b1; \
	doodle_left_alpha[4][75] = 1'b1; \
	doodle_left_alpha[4][76] = 1'b1; \
	doodle_left_alpha[4][77] = 1'b1; \
	doodle_left_alpha[4][78] = 1'b1; \
	doodle_left_alpha[4][79] = 1'b1; \
	doodle_left_alpha[5][0] = 1'b1; \
	doodle_left_alpha[5][1] = 1'b1; \
	doodle_left_alpha[5][2] = 1'b1; \
	doodle_left_alpha[5][3] = 1'b1; \
	doodle_left_alpha[5][4] = 1'b1; \
	doodle_left_alpha[5][5] = 1'b1; \
	doodle_left_alpha[5][6] = 1'b1; \
	doodle_left_alpha[5][7] = 1'b1; \
	doodle_left_alpha[5][8] = 1'b1; \
	doodle_left_alpha[5][9] = 1'b1; \
	doodle_left_alpha[5][10] = 1'b1; \
	doodle_left_alpha[5][11] = 1'b1; \
	doodle_left_alpha[5][12] = 1'b1; \
	doodle_left_alpha[5][13] = 1'b1; \
	doodle_left_alpha[5][14] = 1'b1; \
	doodle_left_alpha[5][15] = 1'b1; \
	doodle_left_alpha[5][16] = 1'b1; \
	doodle_left_alpha[5][17] = 1'b1; \
	doodle_left_alpha[5][18] = 1'b1; \
	doodle_left_alpha[5][19] = 1'b1; \
	doodle_left_alpha[5][20] = 1'b1; \
	doodle_left_alpha[5][21] = 1'b1; \
	doodle_left_alpha[5][22] = 1'b1; \
	doodle_left_alpha[5][23] = 1'b1; \
	doodle_left_alpha[5][24] = 1'b1; \
	doodle_left_alpha[5][25] = 1'b1; \
	doodle_left_alpha[5][26] = 1'b1; \
	doodle_left_alpha[5][27] = 1'b1; \
	doodle_left_alpha[5][28] = 1'b1; \
	doodle_left_alpha[5][29] = 1'b1; \
	doodle_left_alpha[5][30] = 1'b1; \
	doodle_left_alpha[5][31] = 1'b1; \
	doodle_left_alpha[5][32] = 1'b1; \
	doodle_left_alpha[5][33] = 1'b1; \
	doodle_left_alpha[5][34] = 1'b1; \
	doodle_left_alpha[5][35] = 1'b1; \
	doodle_left_alpha[5][36] = 1'b1; \
	doodle_left_alpha[5][37] = 1'b1; \
	doodle_left_alpha[5][38] = 1'b1; \
	doodle_left_alpha[5][39] = 1'b1; \
	doodle_left_alpha[5][40] = 1'b1; \
	doodle_left_alpha[5][41] = 1'b1; \
	doodle_left_alpha[5][42] = 1'b1; \
	doodle_left_alpha[5][43] = 1'b1; \
	doodle_left_alpha[5][44] = 1'b1; \
	doodle_left_alpha[5][45] = 1'b1; \
	doodle_left_alpha[5][46] = 1'b1; \
	doodle_left_alpha[5][47] = 1'b1; \
	doodle_left_alpha[5][48] = 1'b1; \
	doodle_left_alpha[5][49] = 1'b1; \
	doodle_left_alpha[5][50] = 1'b1; \
	doodle_left_alpha[5][51] = 1'b1; \
	doodle_left_alpha[5][52] = 1'b1; \
	doodle_left_alpha[5][53] = 1'b1; \
	doodle_left_alpha[5][54] = 1'b1; \
	doodle_left_alpha[5][55] = 1'b1; \
	doodle_left_alpha[5][56] = 1'b1; \
	doodle_left_alpha[5][57] = 1'b1; \
	doodle_left_alpha[5][58] = 1'b1; \
	doodle_left_alpha[5][59] = 1'b1; \
	doodle_left_alpha[5][60] = 1'b1; \
	doodle_left_alpha[5][61] = 1'b1; \
	doodle_left_alpha[5][62] = 1'b1; \
	doodle_left_alpha[5][63] = 1'b1; \
	doodle_left_alpha[5][64] = 1'b1; \
	doodle_left_alpha[5][65] = 1'b1; \
	doodle_left_alpha[5][66] = 1'b1; \
	doodle_left_alpha[5][67] = 1'b1; \
	doodle_left_alpha[5][68] = 1'b1; \
	doodle_left_alpha[5][69] = 1'b1; \
	doodle_left_alpha[5][70] = 1'b1; \
	doodle_left_alpha[5][71] = 1'b1; \
	doodle_left_alpha[5][72] = 1'b1; \
	doodle_left_alpha[5][73] = 1'b1; \
	doodle_left_alpha[5][74] = 1'b1; \
	doodle_left_alpha[5][75] = 1'b1; \
	doodle_left_alpha[5][76] = 1'b1; \
	doodle_left_alpha[5][77] = 1'b1; \
	doodle_left_alpha[5][78] = 1'b1; \
	doodle_left_alpha[5][79] = 1'b1; \
	doodle_left_alpha[6][0] = 1'b1; \
	doodle_left_alpha[6][1] = 1'b1; \
	doodle_left_alpha[6][2] = 1'b1; \
	doodle_left_alpha[6][3] = 1'b1; \
	doodle_left_alpha[6][4] = 1'b1; \
	doodle_left_alpha[6][5] = 1'b1; \
	doodle_left_alpha[6][6] = 1'b1; \
	doodle_left_alpha[6][7] = 1'b1; \
	doodle_left_alpha[6][8] = 1'b1; \
	doodle_left_alpha[6][9] = 1'b1; \
	doodle_left_alpha[6][10] = 1'b1; \
	doodle_left_alpha[6][11] = 1'b1; \
	doodle_left_alpha[6][12] = 1'b1; \
	doodle_left_alpha[6][13] = 1'b1; \
	doodle_left_alpha[6][14] = 1'b1; \
	doodle_left_alpha[6][15] = 1'b1; \
	doodle_left_alpha[6][16] = 1'b1; \
	doodle_left_alpha[6][17] = 1'b1; \
	doodle_left_alpha[6][18] = 1'b1; \
	doodle_left_alpha[6][19] = 1'b1; \
	doodle_left_alpha[6][20] = 1'b1; \
	doodle_left_alpha[6][21] = 1'b1; \
	doodle_left_alpha[6][22] = 1'b1; \
	doodle_left_alpha[6][23] = 1'b1; \
	doodle_left_alpha[6][24] = 1'b1; \
	doodle_left_alpha[6][25] = 1'b1; \
	doodle_left_alpha[6][26] = 1'b1; \
	doodle_left_alpha[6][27] = 1'b1; \
	doodle_left_alpha[6][28] = 1'b1; \
	doodle_left_alpha[6][29] = 1'b1; \
	doodle_left_alpha[6][30] = 1'b1; \
	doodle_left_alpha[6][31] = 1'b1; \
	doodle_left_alpha[6][32] = 1'b1; \
	doodle_left_alpha[6][33] = 1'b1; \
	doodle_left_alpha[6][34] = 1'b1; \
	doodle_left_alpha[6][35] = 1'b1; \
	doodle_left_alpha[6][36] = 1'b1; \
	doodle_left_alpha[6][37] = 1'b1; \
	doodle_left_alpha[6][38] = 1'b1; \
	doodle_left_alpha[6][39] = 1'b1; \
	doodle_left_alpha[6][40] = 1'b1; \
	doodle_left_alpha[6][41] = 1'b1; \
	doodle_left_alpha[6][42] = 1'b1; \
	doodle_left_alpha[6][43] = 1'b1; \
	doodle_left_alpha[6][44] = 1'b1; \
	doodle_left_alpha[6][45] = 1'b1; \
	doodle_left_alpha[6][46] = 1'b1; \
	doodle_left_alpha[6][47] = 1'b1; \
	doodle_left_alpha[6][48] = 1'b1; \
	doodle_left_alpha[6][49] = 1'b1; \
	doodle_left_alpha[6][50] = 1'b1; \
	doodle_left_alpha[6][51] = 1'b1; \
	doodle_left_alpha[6][52] = 1'b1; \
	doodle_left_alpha[6][53] = 1'b1; \
	doodle_left_alpha[6][54] = 1'b1; \
	doodle_left_alpha[6][55] = 1'b1; \
	doodle_left_alpha[6][56] = 1'b1; \
	doodle_left_alpha[6][57] = 1'b1; \
	doodle_left_alpha[6][58] = 1'b1; \
	doodle_left_alpha[6][59] = 1'b1; \
	doodle_left_alpha[6][60] = 1'b1; \
	doodle_left_alpha[6][61] = 1'b1; \
	doodle_left_alpha[6][62] = 1'b1; \
	doodle_left_alpha[6][63] = 1'b1; \
	doodle_left_alpha[6][64] = 1'b1; \
	doodle_left_alpha[6][65] = 1'b1; \
	doodle_left_alpha[6][66] = 1'b1; \
	doodle_left_alpha[6][67] = 1'b1; \
	doodle_left_alpha[6][68] = 1'b1; \
	doodle_left_alpha[6][69] = 1'b1; \
	doodle_left_alpha[6][70] = 1'b1; \
	doodle_left_alpha[6][71] = 1'b1; \
	doodle_left_alpha[6][72] = 1'b1; \
	doodle_left_alpha[6][73] = 1'b1; \
	doodle_left_alpha[6][74] = 1'b1; \
	doodle_left_alpha[6][75] = 1'b1; \
	doodle_left_alpha[6][76] = 1'b1; \
	doodle_left_alpha[6][77] = 1'b1; \
	doodle_left_alpha[6][78] = 1'b1; \
	doodle_left_alpha[6][79] = 1'b1; \
	doodle_left_alpha[7][0] = 1'b1; \
	doodle_left_alpha[7][1] = 1'b1; \
	doodle_left_alpha[7][2] = 1'b1; \
	doodle_left_alpha[7][3] = 1'b1; \
	doodle_left_alpha[7][4] = 1'b1; \
	doodle_left_alpha[7][5] = 1'b1; \
	doodle_left_alpha[7][6] = 1'b1; \
	doodle_left_alpha[7][7] = 1'b1; \
	doodle_left_alpha[7][8] = 1'b1; \
	doodle_left_alpha[7][9] = 1'b1; \
	doodle_left_alpha[7][10] = 1'b1; \
	doodle_left_alpha[7][11] = 1'b1; \
	doodle_left_alpha[7][12] = 1'b1; \
	doodle_left_alpha[7][13] = 1'b1; \
	doodle_left_alpha[7][14] = 1'b1; \
	doodle_left_alpha[7][15] = 1'b1; \
	doodle_left_alpha[7][16] = 1'b1; \
	doodle_left_alpha[7][17] = 1'b1; \
	doodle_left_alpha[7][18] = 1'b1; \
	doodle_left_alpha[7][19] = 1'b1; \
	doodle_left_alpha[7][20] = 1'b1; \
	doodle_left_alpha[7][21] = 1'b1; \
	doodle_left_alpha[7][22] = 1'b1; \
	doodle_left_alpha[7][23] = 1'b1; \
	doodle_left_alpha[7][24] = 1'b1; \
	doodle_left_alpha[7][25] = 1'b1; \
	doodle_left_alpha[7][26] = 1'b1; \
	doodle_left_alpha[7][27] = 1'b1; \
	doodle_left_alpha[7][28] = 1'b1; \
	doodle_left_alpha[7][29] = 1'b1; \
	doodle_left_alpha[7][30] = 1'b1; \
	doodle_left_alpha[7][31] = 1'b1; \
	doodle_left_alpha[7][32] = 1'b1; \
	doodle_left_alpha[7][33] = 1'b1; \
	doodle_left_alpha[7][34] = 1'b1; \
	doodle_left_alpha[7][35] = 1'b1; \
	doodle_left_alpha[7][36] = 1'b1; \
	doodle_left_alpha[7][37] = 1'b1; \
	doodle_left_alpha[7][38] = 1'b1; \
	doodle_left_alpha[7][39] = 1'b1; \
	doodle_left_alpha[7][40] = 1'b1; \
	doodle_left_alpha[7][41] = 1'b1; \
	doodle_left_alpha[7][42] = 1'b1; \
	doodle_left_alpha[7][43] = 1'b1; \
	doodle_left_alpha[7][44] = 1'b1; \
	doodle_left_alpha[7][45] = 1'b1; \
	doodle_left_alpha[7][46] = 1'b1; \
	doodle_left_alpha[7][47] = 1'b1; \
	doodle_left_alpha[7][48] = 1'b1; \
	doodle_left_alpha[7][49] = 1'b1; \
	doodle_left_alpha[7][50] = 1'b1; \
	doodle_left_alpha[7][51] = 1'b1; \
	doodle_left_alpha[7][52] = 1'b1; \
	doodle_left_alpha[7][53] = 1'b1; \
	doodle_left_alpha[7][54] = 1'b1; \
	doodle_left_alpha[7][55] = 1'b1; \
	doodle_left_alpha[7][56] = 1'b1; \
	doodle_left_alpha[7][57] = 1'b1; \
	doodle_left_alpha[7][58] = 1'b1; \
	doodle_left_alpha[7][59] = 1'b1; \
	doodle_left_alpha[7][60] = 1'b1; \
	doodle_left_alpha[7][61] = 1'b1; \
	doodle_left_alpha[7][62] = 1'b1; \
	doodle_left_alpha[7][63] = 1'b1; \
	doodle_left_alpha[7][64] = 1'b1; \
	doodle_left_alpha[7][65] = 1'b1; \
	doodle_left_alpha[7][66] = 1'b1; \
	doodle_left_alpha[7][67] = 1'b1; \
	doodle_left_alpha[7][68] = 1'b1; \
	doodle_left_alpha[7][69] = 1'b1; \
	doodle_left_alpha[7][70] = 1'b1; \
	doodle_left_alpha[7][71] = 1'b1; \
	doodle_left_alpha[7][72] = 1'b1; \
	doodle_left_alpha[7][73] = 1'b1; \
	doodle_left_alpha[7][74] = 1'b1; \
	doodle_left_alpha[7][75] = 1'b1; \
	doodle_left_alpha[7][76] = 1'b1; \
	doodle_left_alpha[7][77] = 1'b1; \
	doodle_left_alpha[7][78] = 1'b1; \
	doodle_left_alpha[7][79] = 1'b1; \
	doodle_left_alpha[8][0] = 1'b1; \
	doodle_left_alpha[8][1] = 1'b1; \
	doodle_left_alpha[8][2] = 1'b1; \
	doodle_left_alpha[8][3] = 1'b1; \
	doodle_left_alpha[8][4] = 1'b1; \
	doodle_left_alpha[8][5] = 1'b1; \
	doodle_left_alpha[8][6] = 1'b1; \
	doodle_left_alpha[8][7] = 1'b1; \
	doodle_left_alpha[8][8] = 1'b1; \
	doodle_left_alpha[8][9] = 1'b1; \
	doodle_left_alpha[8][10] = 1'b1; \
	doodle_left_alpha[8][11] = 1'b1; \
	doodle_left_alpha[8][12] = 1'b1; \
	doodle_left_alpha[8][13] = 1'b1; \
	doodle_left_alpha[8][14] = 1'b1; \
	doodle_left_alpha[8][15] = 1'b1; \
	doodle_left_alpha[8][16] = 1'b1; \
	doodle_left_alpha[8][17] = 1'b1; \
	doodle_left_alpha[8][18] = 1'b1; \
	doodle_left_alpha[8][19] = 1'b1; \
	doodle_left_alpha[8][20] = 1'b1; \
	doodle_left_alpha[8][21] = 1'b1; \
	doodle_left_alpha[8][22] = 1'b1; \
	doodle_left_alpha[8][23] = 1'b1; \
	doodle_left_alpha[8][24] = 1'b1; \
	doodle_left_alpha[8][25] = 1'b1; \
	doodle_left_alpha[8][26] = 1'b1; \
	doodle_left_alpha[8][27] = 1'b1; \
	doodle_left_alpha[8][28] = 1'b1; \
	doodle_left_alpha[8][29] = 1'b1; \
	doodle_left_alpha[8][30] = 1'b1; \
	doodle_left_alpha[8][31] = 1'b1; \
	doodle_left_alpha[8][32] = 1'b1; \
	doodle_left_alpha[8][33] = 1'b1; \
	doodle_left_alpha[8][34] = 1'b1; \
	doodle_left_alpha[8][35] = 1'b1; \
	doodle_left_alpha[8][36] = 1'b1; \
	doodle_left_alpha[8][37] = 1'b1; \
	doodle_left_alpha[8][38] = 1'b1; \
	doodle_left_alpha[8][39] = 1'b1; \
	doodle_left_alpha[8][40] = 1'b1; \
	doodle_left_alpha[8][41] = 1'b1; \
	doodle_left_alpha[8][42] = 1'b1; \
	doodle_left_alpha[8][43] = 1'b1; \
	doodle_left_alpha[8][44] = 1'b1; \
	doodle_left_alpha[8][45] = 1'b1; \
	doodle_left_alpha[8][46] = 1'b1; \
	doodle_left_alpha[8][47] = 1'b1; \
	doodle_left_alpha[8][48] = 1'b1; \
	doodle_left_alpha[8][49] = 1'b1; \
	doodle_left_alpha[8][50] = 1'b1; \
	doodle_left_alpha[8][51] = 1'b1; \
	doodle_left_alpha[8][52] = 1'b1; \
	doodle_left_alpha[8][53] = 1'b1; \
	doodle_left_alpha[8][54] = 1'b1; \
	doodle_left_alpha[8][55] = 1'b1; \
	doodle_left_alpha[8][56] = 1'b1; \
	doodle_left_alpha[8][57] = 1'b1; \
	doodle_left_alpha[8][58] = 1'b1; \
	doodle_left_alpha[8][59] = 1'b1; \
	doodle_left_alpha[8][60] = 1'b1; \
	doodle_left_alpha[8][61] = 1'b1; \
	doodle_left_alpha[8][62] = 1'b1; \
	doodle_left_alpha[8][63] = 1'b1; \
	doodle_left_alpha[8][64] = 1'b1; \
	doodle_left_alpha[8][65] = 1'b1; \
	doodle_left_alpha[8][66] = 1'b1; \
	doodle_left_alpha[8][67] = 1'b1; \
	doodle_left_alpha[8][68] = 1'b1; \
	doodle_left_alpha[8][69] = 1'b1; \
	doodle_left_alpha[8][70] = 1'b1; \
	doodle_left_alpha[8][71] = 1'b1; \
	doodle_left_alpha[8][72] = 1'b1; \
	doodle_left_alpha[8][73] = 1'b1; \
	doodle_left_alpha[8][74] = 1'b1; \
	doodle_left_alpha[8][75] = 1'b1; \
	doodle_left_alpha[8][76] = 1'b1; \
	doodle_left_alpha[8][77] = 1'b1; \
	doodle_left_alpha[8][78] = 1'b1; \
	doodle_left_alpha[8][79] = 1'b1; \
	doodle_left_alpha[9][0] = 1'b1; \
	doodle_left_alpha[9][1] = 1'b1; \
	doodle_left_alpha[9][2] = 1'b1; \
	doodle_left_alpha[9][3] = 1'b1; \
	doodle_left_alpha[9][4] = 1'b1; \
	doodle_left_alpha[9][5] = 1'b1; \
	doodle_left_alpha[9][6] = 1'b1; \
	doodle_left_alpha[9][7] = 1'b1; \
	doodle_left_alpha[9][8] = 1'b1; \
	doodle_left_alpha[9][9] = 1'b1; \
	doodle_left_alpha[9][10] = 1'b1; \
	doodle_left_alpha[9][11] = 1'b1; \
	doodle_left_alpha[9][12] = 1'b1; \
	doodle_left_alpha[9][13] = 1'b1; \
	doodle_left_alpha[9][14] = 1'b1; \
	doodle_left_alpha[9][15] = 1'b1; \
	doodle_left_alpha[9][16] = 1'b1; \
	doodle_left_alpha[9][17] = 1'b1; \
	doodle_left_alpha[9][18] = 1'b1; \
	doodle_left_alpha[9][19] = 1'b1; \
	doodle_left_alpha[9][20] = 1'b1; \
	doodle_left_alpha[9][21] = 1'b1; \
	doodle_left_alpha[9][22] = 1'b1; \
	doodle_left_alpha[9][23] = 1'b1; \
	doodle_left_alpha[9][24] = 1'b1; \
	doodle_left_alpha[9][25] = 1'b1; \
	doodle_left_alpha[9][26] = 1'b1; \
	doodle_left_alpha[9][27] = 1'b1; \
	doodle_left_alpha[9][28] = 1'b1; \
	doodle_left_alpha[9][29] = 1'b1; \
	doodle_left_alpha[9][30] = 1'b1; \
	doodle_left_alpha[9][31] = 1'b1; \
	doodle_left_alpha[9][32] = 1'b1; \
	doodle_left_alpha[9][33] = 1'b1; \
	doodle_left_alpha[9][34] = 1'b1; \
	doodle_left_alpha[9][35] = 1'b1; \
	doodle_left_alpha[9][36] = 1'b1; \
	doodle_left_alpha[9][37] = 1'b1; \
	doodle_left_alpha[9][38] = 1'b1; \
	doodle_left_alpha[9][39] = 1'b1; \
	doodle_left_alpha[9][40] = 1'b1; \
	doodle_left_alpha[9][41] = 1'b1; \
	doodle_left_alpha[9][42] = 1'b1; \
	doodle_left_alpha[9][43] = 1'b1; \
	doodle_left_alpha[9][44] = 1'b1; \
	doodle_left_alpha[9][45] = 1'b1; \
	doodle_left_alpha[9][46] = 1'b1; \
	doodle_left_alpha[9][47] = 1'b1; \
	doodle_left_alpha[9][48] = 1'b1; \
	doodle_left_alpha[9][49] = 1'b1; \
	doodle_left_alpha[9][50] = 1'b1; \
	doodle_left_alpha[9][51] = 1'b1; \
	doodle_left_alpha[9][52] = 1'b1; \
	doodle_left_alpha[9][53] = 1'b1; \
	doodle_left_alpha[9][54] = 1'b1; \
	doodle_left_alpha[9][55] = 1'b1; \
	doodle_left_alpha[9][56] = 1'b1; \
	doodle_left_alpha[9][57] = 1'b1; \
	doodle_left_alpha[9][58] = 1'b1; \
	doodle_left_alpha[9][59] = 1'b1; \
	doodle_left_alpha[9][60] = 1'b1; \
	doodle_left_alpha[9][61] = 1'b1; \
	doodle_left_alpha[9][62] = 1'b1; \
	doodle_left_alpha[9][63] = 1'b1; \
	doodle_left_alpha[9][64] = 1'b1; \
	doodle_left_alpha[9][65] = 1'b1; \
	doodle_left_alpha[9][66] = 1'b1; \
	doodle_left_alpha[9][67] = 1'b1; \
	doodle_left_alpha[9][68] = 1'b1; \
	doodle_left_alpha[9][69] = 1'b1; \
	doodle_left_alpha[9][70] = 1'b1; \
	doodle_left_alpha[9][71] = 1'b1; \
	doodle_left_alpha[9][72] = 1'b1; \
	doodle_left_alpha[9][73] = 1'b1; \
	doodle_left_alpha[9][74] = 1'b1; \
	doodle_left_alpha[9][75] = 1'b1; \
	doodle_left_alpha[9][76] = 1'b1; \
	doodle_left_alpha[9][77] = 1'b1; \
	doodle_left_alpha[9][78] = 1'b1; \
	doodle_left_alpha[9][79] = 1'b1; \
	doodle_left_alpha[10][0] = 1'b1; \
	doodle_left_alpha[10][1] = 1'b1; \
	doodle_left_alpha[10][2] = 1'b1; \
	doodle_left_alpha[10][3] = 1'b1; \
	doodle_left_alpha[10][4] = 1'b1; \
	doodle_left_alpha[10][5] = 1'b1; \
	doodle_left_alpha[10][6] = 1'b1; \
	doodle_left_alpha[10][7] = 1'b1; \
	doodle_left_alpha[10][8] = 1'b1; \
	doodle_left_alpha[10][9] = 1'b1; \
	doodle_left_alpha[10][10] = 1'b1; \
	doodle_left_alpha[10][11] = 1'b1; \
	doodle_left_alpha[10][12] = 1'b1; \
	doodle_left_alpha[10][13] = 1'b1; \
	doodle_left_alpha[10][14] = 1'b1; \
	doodle_left_alpha[10][15] = 1'b1; \
	doodle_left_alpha[10][16] = 1'b1; \
	doodle_left_alpha[10][17] = 1'b1; \
	doodle_left_alpha[10][18] = 1'b1; \
	doodle_left_alpha[10][19] = 1'b1; \
	doodle_left_alpha[10][20] = 1'b1; \
	doodle_left_alpha[10][21] = 1'b1; \
	doodle_left_alpha[10][22] = 1'b1; \
	doodle_left_alpha[10][23] = 1'b1; \
	doodle_left_alpha[10][24] = 1'b1; \
	doodle_left_alpha[10][25] = 1'b1; \
	doodle_left_alpha[10][26] = 1'b1; \
	doodle_left_alpha[10][27] = 1'b1; \
	doodle_left_alpha[10][28] = 1'b1; \
	doodle_left_alpha[10][29] = 1'b1; \
	doodle_left_alpha[10][30] = 1'b1; \
	doodle_left_alpha[10][31] = 1'b1; \
	doodle_left_alpha[10][32] = 1'b1; \
	doodle_left_alpha[10][33] = 1'b1; \
	doodle_left_alpha[10][34] = 1'b1; \
	doodle_left_alpha[10][35] = 1'b1; \
	doodle_left_alpha[10][36] = 1'b1; \
	doodle_left_alpha[10][37] = 1'b1; \
	doodle_left_alpha[10][38] = 1'b1; \
	doodle_left_alpha[10][39] = 1'b1; \
	doodle_left_alpha[10][40] = 1'b1; \
	doodle_left_alpha[10][41] = 1'b1; \
	doodle_left_alpha[10][42] = 1'b1; \
	doodle_left_alpha[10][43] = 1'b1; \
	doodle_left_alpha[10][44] = 1'b1; \
	doodle_left_alpha[10][45] = 1'b1; \
	doodle_left_alpha[10][46] = 1'b1; \
	doodle_left_alpha[10][47] = 1'b1; \
	doodle_left_alpha[10][48] = 1'b1; \
	doodle_left_alpha[10][49] = 1'b1; \
	doodle_left_alpha[10][50] = 1'b1; \
	doodle_left_alpha[10][51] = 1'b1; \
	doodle_left_alpha[10][52] = 1'b1; \
	doodle_left_alpha[10][53] = 1'b1; \
	doodle_left_alpha[10][54] = 1'b1; \
	doodle_left_alpha[10][55] = 1'b1; \
	doodle_left_alpha[10][56] = 1'b1; \
	doodle_left_alpha[10][57] = 1'b1; \
	doodle_left_alpha[10][58] = 1'b1; \
	doodle_left_alpha[10][59] = 1'b1; \
	doodle_left_alpha[10][60] = 1'b1; \
	doodle_left_alpha[10][61] = 1'b1; \
	doodle_left_alpha[10][62] = 1'b1; \
	doodle_left_alpha[10][63] = 1'b1; \
	doodle_left_alpha[10][64] = 1'b1; \
	doodle_left_alpha[10][65] = 1'b1; \
	doodle_left_alpha[10][66] = 1'b1; \
	doodle_left_alpha[10][67] = 1'b1; \
	doodle_left_alpha[10][68] = 1'b1; \
	doodle_left_alpha[10][69] = 1'b1; \
	doodle_left_alpha[10][70] = 1'b1; \
	doodle_left_alpha[10][71] = 1'b1; \
	doodle_left_alpha[10][72] = 1'b1; \
	doodle_left_alpha[10][73] = 1'b1; \
	doodle_left_alpha[10][74] = 1'b1; \
	doodle_left_alpha[10][75] = 1'b1; \
	doodle_left_alpha[10][76] = 1'b1; \
	doodle_left_alpha[10][77] = 1'b1; \
	doodle_left_alpha[10][78] = 1'b1; \
	doodle_left_alpha[10][79] = 1'b1; \
	doodle_left_alpha[11][0] = 1'b1; \
	doodle_left_alpha[11][1] = 1'b1; \
	doodle_left_alpha[11][2] = 1'b1; \
	doodle_left_alpha[11][3] = 1'b1; \
	doodle_left_alpha[11][4] = 1'b1; \
	doodle_left_alpha[11][5] = 1'b1; \
	doodle_left_alpha[11][6] = 1'b1; \
	doodle_left_alpha[11][7] = 1'b1; \
	doodle_left_alpha[11][8] = 1'b1; \
	doodle_left_alpha[11][9] = 1'b1; \
	doodle_left_alpha[11][10] = 1'b1; \
	doodle_left_alpha[11][11] = 1'b1; \
	doodle_left_alpha[11][12] = 1'b1; \
	doodle_left_alpha[11][13] = 1'b1; \
	doodle_left_alpha[11][14] = 1'b1; \
	doodle_left_alpha[11][15] = 1'b1; \
	doodle_left_alpha[11][16] = 1'b1; \
	doodle_left_alpha[11][17] = 1'b1; \
	doodle_left_alpha[11][18] = 1'b1; \
	doodle_left_alpha[11][19] = 1'b1; \
	doodle_left_alpha[11][20] = 1'b1; \
	doodle_left_alpha[11][21] = 1'b1; \
	doodle_left_alpha[11][22] = 1'b1; \
	doodle_left_alpha[11][23] = 1'b1; \
	doodle_left_alpha[11][24] = 1'b1; \
	doodle_left_alpha[11][25] = 1'b1; \
	doodle_left_alpha[11][26] = 1'b1; \
	doodle_left_alpha[11][27] = 1'b1; \
	doodle_left_alpha[11][28] = 1'b1; \
	doodle_left_alpha[11][29] = 1'b1; \
	doodle_left_alpha[11][30] = 1'b1; \
	doodle_left_alpha[11][31] = 1'b1; \
	doodle_left_alpha[11][32] = 1'b1; \
	doodle_left_alpha[11][33] = 1'b1; \
	doodle_left_alpha[11][34] = 1'b1; \
	doodle_left_alpha[11][35] = 1'b1; \
	doodle_left_alpha[11][36] = 1'b1; \
	doodle_left_alpha[11][37] = 1'b1; \
	doodle_left_alpha[11][38] = 1'b1; \
	doodle_left_alpha[11][39] = 1'b1; \
	doodle_left_alpha[11][40] = 1'b1; \
	doodle_left_alpha[11][41] = 1'b1; \
	doodle_left_alpha[11][42] = 1'b1; \
	doodle_left_alpha[11][43] = 1'b1; \
	doodle_left_alpha[11][44] = 1'b1; \
	doodle_left_alpha[11][45] = 1'b1; \
	doodle_left_alpha[11][46] = 1'b1; \
	doodle_left_alpha[11][47] = 1'b1; \
	doodle_left_alpha[11][48] = 1'b1; \
	doodle_left_alpha[11][49] = 1'b1; \
	doodle_left_alpha[11][50] = 1'b1; \
	doodle_left_alpha[11][51] = 1'b1; \
	doodle_left_alpha[11][52] = 1'b1; \
	doodle_left_alpha[11][53] = 1'b1; \
	doodle_left_alpha[11][54] = 1'b1; \
	doodle_left_alpha[11][55] = 1'b1; \
	doodle_left_alpha[11][56] = 1'b1; \
	doodle_left_alpha[11][57] = 1'b1; \
	doodle_left_alpha[11][58] = 1'b1; \
	doodle_left_alpha[11][59] = 1'b1; \
	doodle_left_alpha[11][60] = 1'b1; \
	doodle_left_alpha[11][61] = 1'b1; \
	doodle_left_alpha[11][62] = 1'b1; \
	doodle_left_alpha[11][63] = 1'b1; \
	doodle_left_alpha[11][64] = 1'b1; \
	doodle_left_alpha[11][65] = 1'b1; \
	doodle_left_alpha[11][66] = 1'b1; \
	doodle_left_alpha[11][67] = 1'b1; \
	doodle_left_alpha[11][68] = 1'b1; \
	doodle_left_alpha[11][69] = 1'b1; \
	doodle_left_alpha[11][70] = 1'b1; \
	doodle_left_alpha[11][71] = 1'b1; \
	doodle_left_alpha[11][72] = 1'b1; \
	doodle_left_alpha[11][73] = 1'b1; \
	doodle_left_alpha[11][74] = 1'b1; \
	doodle_left_alpha[11][75] = 1'b1; \
	doodle_left_alpha[11][76] = 1'b1; \
	doodle_left_alpha[11][77] = 1'b1; \
	doodle_left_alpha[11][78] = 1'b1; \
	doodle_left_alpha[11][79] = 1'b1; \
	doodle_left_alpha[12][0] = 1'b1; \
	doodle_left_alpha[12][1] = 1'b1; \
	doodle_left_alpha[12][2] = 1'b1; \
	doodle_left_alpha[12][3] = 1'b1; \
	doodle_left_alpha[12][4] = 1'b1; \
	doodle_left_alpha[12][5] = 1'b1; \
	doodle_left_alpha[12][6] = 1'b1; \
	doodle_left_alpha[12][7] = 1'b1; \
	doodle_left_alpha[12][8] = 1'b1; \
	doodle_left_alpha[12][9] = 1'b1; \
	doodle_left_alpha[12][10] = 1'b1; \
	doodle_left_alpha[12][11] = 1'b1; \
	doodle_left_alpha[12][12] = 1'b1; \
	doodle_left_alpha[12][13] = 1'b1; \
	doodle_left_alpha[12][14] = 1'b1; \
	doodle_left_alpha[12][15] = 1'b1; \
	doodle_left_alpha[12][16] = 1'b1; \
	doodle_left_alpha[12][17] = 1'b1; \
	doodle_left_alpha[12][18] = 1'b1; \
	doodle_left_alpha[12][19] = 1'b1; \
	doodle_left_alpha[12][20] = 1'b1; \
	doodle_left_alpha[12][21] = 1'b1; \
	doodle_left_alpha[12][22] = 1'b1; \
	doodle_left_alpha[12][23] = 1'b1; \
	doodle_left_alpha[12][24] = 1'b1; \
	doodle_left_alpha[12][25] = 1'b1; \
	doodle_left_alpha[12][26] = 1'b1; \
	doodle_left_alpha[12][27] = 1'b1; \
	doodle_left_alpha[12][28] = 1'b1; \
	doodle_left_alpha[12][29] = 1'b1; \
	doodle_left_alpha[12][30] = 1'b1; \
	doodle_left_alpha[12][31] = 1'b1; \
	doodle_left_alpha[12][32] = 1'b1; \
	doodle_left_alpha[12][33] = 1'b1; \
	doodle_left_alpha[12][34] = 1'b1; \
	doodle_left_alpha[12][35] = 1'b1; \
	doodle_left_alpha[12][36] = 1'b1; \
	doodle_left_alpha[12][37] = 1'b1; \
	doodle_left_alpha[12][38] = 1'b1; \
	doodle_left_alpha[12][39] = 1'b1; \
	doodle_left_alpha[12][40] = 1'b1; \
	doodle_left_alpha[12][41] = 1'b1; \
	doodle_left_alpha[12][42] = 1'b1; \
	doodle_left_alpha[12][43] = 1'b1; \
	doodle_left_alpha[12][44] = 1'b1; \
	doodle_left_alpha[12][45] = 1'b1; \
	doodle_left_alpha[12][46] = 1'b1; \
	doodle_left_alpha[12][47] = 1'b1; \
	doodle_left_alpha[12][48] = 1'b1; \
	doodle_left_alpha[12][49] = 1'b1; \
	doodle_left_alpha[12][50] = 1'b1; \
	doodle_left_alpha[12][51] = 1'b1; \
	doodle_left_alpha[12][52] = 1'b1; \
	doodle_left_alpha[12][53] = 1'b1; \
	doodle_left_alpha[12][54] = 1'b1; \
	doodle_left_alpha[12][55] = 1'b1; \
	doodle_left_alpha[12][56] = 1'b1; \
	doodle_left_alpha[12][57] = 1'b1; \
	doodle_left_alpha[12][58] = 1'b1; \
	doodle_left_alpha[12][59] = 1'b1; \
	doodle_left_alpha[12][60] = 1'b1; \
	doodle_left_alpha[12][61] = 1'b1; \
	doodle_left_alpha[12][62] = 1'b1; \
	doodle_left_alpha[12][63] = 1'b1; \
	doodle_left_alpha[12][64] = 1'b1; \
	doodle_left_alpha[12][65] = 1'b1; \
	doodle_left_alpha[12][66] = 1'b1; \
	doodle_left_alpha[12][67] = 1'b1; \
	doodle_left_alpha[12][68] = 1'b1; \
	doodle_left_alpha[12][69] = 1'b1; \
	doodle_left_alpha[12][70] = 1'b1; \
	doodle_left_alpha[12][71] = 1'b1; \
	doodle_left_alpha[12][72] = 1'b1; \
	doodle_left_alpha[12][73] = 1'b1; \
	doodle_left_alpha[12][74] = 1'b1; \
	doodle_left_alpha[12][75] = 1'b1; \
	doodle_left_alpha[12][76] = 1'b1; \
	doodle_left_alpha[12][77] = 1'b1; \
	doodle_left_alpha[12][78] = 1'b1; \
	doodle_left_alpha[12][79] = 1'b1; \
	doodle_left_alpha[13][0] = 1'b1; \
	doodle_left_alpha[13][1] = 1'b1; \
	doodle_left_alpha[13][2] = 1'b1; \
	doodle_left_alpha[13][3] = 1'b1; \
	doodle_left_alpha[13][4] = 1'b1; \
	doodle_left_alpha[13][5] = 1'b1; \
	doodle_left_alpha[13][6] = 1'b1; \
	doodle_left_alpha[13][7] = 1'b1; \
	doodle_left_alpha[13][8] = 1'b1; \
	doodle_left_alpha[13][9] = 1'b1; \
	doodle_left_alpha[13][10] = 1'b1; \
	doodle_left_alpha[13][11] = 1'b1; \
	doodle_left_alpha[13][12] = 1'b1; \
	doodle_left_alpha[13][13] = 1'b1; \
	doodle_left_alpha[13][14] = 1'b1; \
	doodle_left_alpha[13][15] = 1'b1; \
	doodle_left_alpha[13][16] = 1'b1; \
	doodle_left_alpha[13][17] = 1'b1; \
	doodle_left_alpha[13][18] = 1'b1; \
	doodle_left_alpha[13][19] = 1'b1; \
	doodle_left_alpha[13][20] = 1'b1; \
	doodle_left_alpha[13][21] = 1'b1; \
	doodle_left_alpha[13][22] = 1'b1; \
	doodle_left_alpha[13][23] = 1'b1; \
	doodle_left_alpha[13][24] = 1'b1; \
	doodle_left_alpha[13][25] = 1'b1; \
	doodle_left_alpha[13][26] = 1'b1; \
	doodle_left_alpha[13][27] = 1'b1; \
	doodle_left_alpha[13][28] = 1'b1; \
	doodle_left_alpha[13][29] = 1'b1; \
	doodle_left_alpha[13][30] = 1'b1; \
	doodle_left_alpha[13][31] = 1'b1; \
	doodle_left_alpha[13][32] = 1'b1; \
	doodle_left_alpha[13][33] = 1'b1; \
	doodle_left_alpha[13][34] = 1'b1; \
	doodle_left_alpha[13][35] = 1'b1; \
	doodle_left_alpha[13][36] = 1'b1; \
	doodle_left_alpha[13][37] = 1'b1; \
	doodle_left_alpha[13][38] = 1'b1; \
	doodle_left_alpha[13][39] = 1'b1; \
	doodle_left_alpha[13][40] = 1'b1; \
	doodle_left_alpha[13][41] = 1'b1; \
	doodle_left_alpha[13][42] = 1'b1; \
	doodle_left_alpha[13][43] = 1'b1; \
	doodle_left_alpha[13][44] = 1'b1; \
	doodle_left_alpha[13][45] = 1'b1; \
	doodle_left_alpha[13][46] = 1'b1; \
	doodle_left_alpha[13][47] = 1'b1; \
	doodle_left_alpha[13][48] = 1'b1; \
	doodle_left_alpha[13][49] = 1'b1; \
	doodle_left_alpha[13][50] = 1'b1; \
	doodle_left_alpha[13][51] = 1'b1; \
	doodle_left_alpha[13][52] = 1'b1; \
	doodle_left_alpha[13][53] = 1'b1; \
	doodle_left_alpha[13][54] = 1'b1; \
	doodle_left_alpha[13][55] = 1'b1; \
	doodle_left_alpha[13][56] = 1'b1; \
	doodle_left_alpha[13][57] = 1'b1; \
	doodle_left_alpha[13][58] = 1'b1; \
	doodle_left_alpha[13][59] = 1'b1; \
	doodle_left_alpha[13][60] = 1'b1; \
	doodle_left_alpha[13][61] = 1'b1; \
	doodle_left_alpha[13][62] = 1'b1; \
	doodle_left_alpha[13][63] = 1'b1; \
	doodle_left_alpha[13][64] = 1'b1; \
	doodle_left_alpha[13][65] = 1'b1; \
	doodle_left_alpha[13][66] = 1'b1; \
	doodle_left_alpha[13][67] = 1'b1; \
	doodle_left_alpha[13][68] = 1'b1; \
	doodle_left_alpha[13][69] = 1'b1; \
	doodle_left_alpha[13][70] = 1'b1; \
	doodle_left_alpha[13][71] = 1'b1; \
	doodle_left_alpha[13][72] = 1'b1; \
	doodle_left_alpha[13][73] = 1'b1; \
	doodle_left_alpha[13][74] = 1'b1; \
	doodle_left_alpha[13][75] = 1'b1; \
	doodle_left_alpha[13][76] = 1'b1; \
	doodle_left_alpha[13][77] = 1'b1; \
	doodle_left_alpha[13][78] = 1'b1; \
	doodle_left_alpha[13][79] = 1'b1; \
	doodle_left_alpha[14][0] = 1'b1; \
	doodle_left_alpha[14][1] = 1'b1; \
	doodle_left_alpha[14][2] = 1'b1; \
	doodle_left_alpha[14][3] = 1'b1; \
	doodle_left_alpha[14][4] = 1'b1; \
	doodle_left_alpha[14][5] = 1'b1; \
	doodle_left_alpha[14][6] = 1'b1; \
	doodle_left_alpha[14][7] = 1'b1; \
	doodle_left_alpha[14][8] = 1'b1; \
	doodle_left_alpha[14][9] = 1'b1; \
	doodle_left_alpha[14][10] = 1'b1; \
	doodle_left_alpha[14][11] = 1'b1; \
	doodle_left_alpha[14][12] = 1'b1; \
	doodle_left_alpha[14][13] = 1'b1; \
	doodle_left_alpha[14][14] = 1'b1; \
	doodle_left_alpha[14][15] = 1'b1; \
	doodle_left_alpha[14][16] = 1'b1; \
	doodle_left_alpha[14][17] = 1'b1; \
	doodle_left_alpha[14][18] = 1'b1; \
	doodle_left_alpha[14][19] = 1'b1; \
	doodle_left_alpha[14][20] = 1'b1; \
	doodle_left_alpha[14][21] = 1'b1; \
	doodle_left_alpha[14][22] = 1'b1; \
	doodle_left_alpha[14][23] = 1'b1; \
	doodle_left_alpha[14][24] = 1'b1; \
	doodle_left_alpha[14][25] = 1'b1; \
	doodle_left_alpha[14][26] = 1'b1; \
	doodle_left_alpha[14][27] = 1'b1; \
	doodle_left_alpha[14][28] = 1'b1; \
	doodle_left_alpha[14][29] = 1'b1; \
	doodle_left_alpha[14][30] = 1'b1; \
	doodle_left_alpha[14][31] = 1'b1; \
	doodle_left_alpha[14][32] = 1'b1; \
	doodle_left_alpha[14][33] = 1'b1; \
	doodle_left_alpha[14][34] = 1'b1; \
	doodle_left_alpha[14][35] = 1'b1; \
	doodle_left_alpha[14][36] = 1'b1; \
	doodle_left_alpha[14][37] = 1'b1; \
	doodle_left_alpha[14][38] = 1'b1; \
	doodle_left_alpha[14][39] = 1'b1; \
	doodle_left_alpha[14][40] = 1'b1; \
	doodle_left_alpha[14][41] = 1'b1; \
	doodle_left_alpha[14][42] = 1'b1; \
	doodle_left_alpha[14][43] = 1'b1; \
	doodle_left_alpha[14][44] = 1'b1; \
	doodle_left_alpha[14][45] = 1'b1; \
	doodle_left_alpha[14][46] = 1'b1; \
	doodle_left_alpha[14][47] = 1'b1; \
	doodle_left_alpha[14][48] = 1'b1; \
	doodle_left_alpha[14][49] = 1'b1; \
	doodle_left_alpha[14][50] = 1'b1; \
	doodle_left_alpha[14][51] = 1'b1; \
	doodle_left_alpha[14][52] = 1'b1; \
	doodle_left_alpha[14][53] = 1'b1; \
	doodle_left_alpha[14][54] = 1'b1; \
	doodle_left_alpha[14][55] = 1'b1; \
	doodle_left_alpha[14][56] = 1'b1; \
	doodle_left_alpha[14][57] = 1'b1; \
	doodle_left_alpha[14][58] = 1'b1; \
	doodle_left_alpha[14][59] = 1'b1; \
	doodle_left_alpha[14][60] = 1'b1; \
	doodle_left_alpha[14][61] = 1'b1; \
	doodle_left_alpha[14][62] = 1'b1; \
	doodle_left_alpha[14][63] = 1'b1; \
	doodle_left_alpha[14][64] = 1'b1; \
	doodle_left_alpha[14][65] = 1'b1; \
	doodle_left_alpha[14][66] = 1'b1; \
	doodle_left_alpha[14][67] = 1'b1; \
	doodle_left_alpha[14][68] = 1'b1; \
	doodle_left_alpha[14][69] = 1'b1; \
	doodle_left_alpha[14][70] = 1'b1; \
	doodle_left_alpha[14][71] = 1'b1; \
	doodle_left_alpha[14][72] = 1'b1; \
	doodle_left_alpha[14][73] = 1'b1; \
	doodle_left_alpha[14][74] = 1'b1; \
	doodle_left_alpha[14][75] = 1'b1; \
	doodle_left_alpha[14][76] = 1'b1; \
	doodle_left_alpha[14][77] = 1'b1; \
	doodle_left_alpha[14][78] = 1'b1; \
	doodle_left_alpha[14][79] = 1'b1; \
	doodle_left_alpha[15][0] = 1'b1; \
	doodle_left_alpha[15][1] = 1'b1; \
	doodle_left_alpha[15][2] = 1'b1; \
	doodle_left_alpha[15][3] = 1'b1; \
	doodle_left_alpha[15][4] = 1'b1; \
	doodle_left_alpha[15][5] = 1'b1; \
	doodle_left_alpha[15][6] = 1'b1; \
	doodle_left_alpha[15][7] = 1'b1; \
	doodle_left_alpha[15][8] = 1'b1; \
	doodle_left_alpha[15][9] = 1'b1; \
	doodle_left_alpha[15][10] = 1'b1; \
	doodle_left_alpha[15][11] = 1'b1; \
	doodle_left_alpha[15][12] = 1'b1; \
	doodle_left_alpha[15][13] = 1'b1; \
	doodle_left_alpha[15][14] = 1'b1; \
	doodle_left_alpha[15][15] = 1'b1; \
	doodle_left_alpha[15][16] = 1'b1; \
	doodle_left_alpha[15][17] = 1'b1; \
	doodle_left_alpha[15][18] = 1'b1; \
	doodle_left_alpha[15][19] = 1'b1; \
	doodle_left_alpha[15][20] = 1'b1; \
	doodle_left_alpha[15][21] = 1'b1; \
	doodle_left_alpha[15][22] = 1'b1; \
	doodle_left_alpha[15][23] = 1'b1; \
	doodle_left_alpha[15][24] = 1'b1; \
	doodle_left_alpha[15][25] = 1'b1; \
	doodle_left_alpha[15][26] = 1'b1; \
	doodle_left_alpha[15][27] = 1'b1; \
	doodle_left_alpha[15][28] = 1'b1; \
	doodle_left_alpha[15][29] = 1'b1; \
	doodle_left_alpha[15][30] = 1'b1; \
	doodle_left_alpha[15][31] = 1'b1; \
	doodle_left_alpha[15][32] = 1'b1; \
	doodle_left_alpha[15][33] = 1'b1; \
	doodle_left_alpha[15][34] = 1'b1; \
	doodle_left_alpha[15][35] = 1'b1; \
	doodle_left_alpha[15][36] = 1'b1; \
	doodle_left_alpha[15][37] = 1'b1; \
	doodle_left_alpha[15][38] = 1'b1; \
	doodle_left_alpha[15][39] = 1'b1; \
	doodle_left_alpha[15][40] = 1'b1; \
	doodle_left_alpha[15][41] = 1'b1; \
	doodle_left_alpha[15][42] = 1'b1; \
	doodle_left_alpha[15][43] = 1'b1; \
	doodle_left_alpha[15][44] = 1'b1; \
	doodle_left_alpha[15][45] = 1'b1; \
	doodle_left_alpha[15][46] = 1'b1; \
	doodle_left_alpha[15][47] = 1'b1; \
	doodle_left_alpha[15][48] = 1'b1; \
	doodle_left_alpha[15][49] = 1'b1; \
	doodle_left_alpha[15][50] = 1'b1; \
	doodle_left_alpha[15][51] = 1'b1; \
	doodle_left_alpha[15][52] = 1'b1; \
	doodle_left_alpha[15][53] = 1'b1; \
	doodle_left_alpha[15][54] = 1'b1; \
	doodle_left_alpha[15][55] = 1'b1; \
	doodle_left_alpha[15][56] = 1'b1; \
	doodle_left_alpha[15][57] = 1'b1; \
	doodle_left_alpha[15][58] = 1'b1; \
	doodle_left_alpha[15][59] = 1'b1; \
	doodle_left_alpha[15][60] = 1'b1; \
	doodle_left_alpha[15][61] = 1'b1; \
	doodle_left_alpha[15][62] = 1'b1; \
	doodle_left_alpha[15][63] = 1'b1; \
	doodle_left_alpha[15][64] = 1'b1; \
	doodle_left_alpha[15][65] = 1'b1; \
	doodle_left_alpha[15][66] = 1'b1; \
	doodle_left_alpha[15][67] = 1'b1; \
	doodle_left_alpha[15][68] = 1'b1; \
	doodle_left_alpha[15][69] = 1'b1; \
	doodle_left_alpha[15][70] = 1'b1; \
	doodle_left_alpha[15][71] = 1'b1; \
	doodle_left_alpha[15][72] = 1'b1; \
	doodle_left_alpha[15][73] = 1'b1; \
	doodle_left_alpha[15][74] = 1'b1; \
	doodle_left_alpha[15][75] = 1'b1; \
	doodle_left_alpha[15][76] = 1'b1; \
	doodle_left_alpha[15][77] = 1'b1; \
	doodle_left_alpha[15][78] = 1'b1; \
	doodle_left_alpha[15][79] = 1'b1; \
	doodle_left_alpha[16][0] = 1'b1; \
	doodle_left_alpha[16][1] = 1'b1; \
	doodle_left_alpha[16][2] = 1'b1; \
	doodle_left_alpha[16][3] = 1'b1; \
	doodle_left_alpha[16][4] = 1'b1; \
	doodle_left_alpha[16][5] = 1'b1; \
	doodle_left_alpha[16][6] = 1'b1; \
	doodle_left_alpha[16][7] = 1'b1; \
	doodle_left_alpha[16][8] = 1'b1; \
	doodle_left_alpha[16][9] = 1'b1; \
	doodle_left_alpha[16][10] = 1'b1; \
	doodle_left_alpha[16][11] = 1'b1; \
	doodle_left_alpha[16][12] = 1'b1; \
	doodle_left_alpha[16][13] = 1'b1; \
	doodle_left_alpha[16][14] = 1'b1; \
	doodle_left_alpha[16][15] = 1'b1; \
	doodle_left_alpha[16][16] = 1'b1; \
	doodle_left_alpha[16][17] = 1'b1; \
	doodle_left_alpha[16][18] = 1'b1; \
	doodle_left_alpha[16][19] = 1'b1; \
	doodle_left_alpha[16][20] = 1'b1; \
	doodle_left_alpha[16][21] = 1'b1; \
	doodle_left_alpha[16][22] = 1'b1; \
	doodle_left_alpha[16][23] = 1'b1; \
	doodle_left_alpha[16][24] = 1'b1; \
	doodle_left_alpha[16][25] = 1'b1; \
	doodle_left_alpha[16][26] = 1'b1; \
	doodle_left_alpha[16][27] = 1'b1; \
	doodle_left_alpha[16][28] = 1'b1; \
	doodle_left_alpha[16][29] = 1'b1; \
	doodle_left_alpha[16][30] = 1'b1; \
	doodle_left_alpha[16][31] = 1'b0; \
	doodle_left_alpha[16][32] = 1'b0; \
	doodle_left_alpha[16][33] = 1'b0; \
	doodle_left_alpha[16][34] = 1'b0; \
	doodle_left_alpha[16][35] = 1'b0; \
	doodle_left_alpha[16][36] = 1'b0; \
	doodle_left_alpha[16][37] = 1'b0; \
	doodle_left_alpha[16][38] = 1'b0; \
	doodle_left_alpha[16][39] = 1'b0; \
	doodle_left_alpha[16][40] = 1'b0; \
	doodle_left_alpha[16][41] = 1'b0; \
	doodle_left_alpha[16][42] = 1'b0; \
	doodle_left_alpha[16][43] = 1'b0; \
	doodle_left_alpha[16][44] = 1'b0; \
	doodle_left_alpha[16][45] = 1'b0; \
	doodle_left_alpha[16][46] = 1'b0; \
	doodle_left_alpha[16][47] = 1'b0; \
	doodle_left_alpha[16][48] = 1'b0; \
	doodle_left_alpha[16][49] = 1'b0; \
	doodle_left_alpha[16][50] = 1'b0; \
	doodle_left_alpha[16][51] = 1'b0; \
	doodle_left_alpha[16][52] = 1'b0; \
	doodle_left_alpha[16][53] = 1'b0; \
	doodle_left_alpha[16][54] = 1'b0; \
	doodle_left_alpha[16][55] = 1'b0; \
	doodle_left_alpha[16][56] = 1'b0; \
	doodle_left_alpha[16][57] = 1'b1; \
	doodle_left_alpha[16][58] = 1'b1; \
	doodle_left_alpha[16][59] = 1'b1; \
	doodle_left_alpha[16][60] = 1'b1; \
	doodle_left_alpha[16][61] = 1'b1; \
	doodle_left_alpha[16][62] = 1'b1; \
	doodle_left_alpha[16][63] = 1'b1; \
	doodle_left_alpha[16][64] = 1'b1; \
	doodle_left_alpha[16][65] = 1'b1; \
	doodle_left_alpha[16][66] = 1'b1; \
	doodle_left_alpha[16][67] = 1'b1; \
	doodle_left_alpha[16][68] = 1'b1; \
	doodle_left_alpha[16][69] = 1'b1; \
	doodle_left_alpha[16][70] = 1'b1; \
	doodle_left_alpha[16][71] = 1'b1; \
	doodle_left_alpha[16][72] = 1'b1; \
	doodle_left_alpha[16][73] = 1'b1; \
	doodle_left_alpha[16][74] = 1'b1; \
	doodle_left_alpha[16][75] = 1'b1; \
	doodle_left_alpha[16][76] = 1'b1; \
	doodle_left_alpha[16][77] = 1'b1; \
	doodle_left_alpha[16][78] = 1'b1; \
	doodle_left_alpha[16][79] = 1'b1; \
	doodle_left_alpha[17][0] = 1'b1; \
	doodle_left_alpha[17][1] = 1'b1; \
	doodle_left_alpha[17][2] = 1'b1; \
	doodle_left_alpha[17][3] = 1'b1; \
	doodle_left_alpha[17][4] = 1'b1; \
	doodle_left_alpha[17][5] = 1'b1; \
	doodle_left_alpha[17][6] = 1'b1; \
	doodle_left_alpha[17][7] = 1'b1; \
	doodle_left_alpha[17][8] = 1'b1; \
	doodle_left_alpha[17][9] = 1'b1; \
	doodle_left_alpha[17][10] = 1'b1; \
	doodle_left_alpha[17][11] = 1'b1; \
	doodle_left_alpha[17][12] = 1'b1; \
	doodle_left_alpha[17][13] = 1'b1; \
	doodle_left_alpha[17][14] = 1'b1; \
	doodle_left_alpha[17][15] = 1'b1; \
	doodle_left_alpha[17][16] = 1'b1; \
	doodle_left_alpha[17][17] = 1'b1; \
	doodle_left_alpha[17][18] = 1'b1; \
	doodle_left_alpha[17][19] = 1'b1; \
	doodle_left_alpha[17][20] = 1'b1; \
	doodle_left_alpha[17][21] = 1'b1; \
	doodle_left_alpha[17][22] = 1'b1; \
	doodle_left_alpha[17][23] = 1'b1; \
	doodle_left_alpha[17][24] = 1'b1; \
	doodle_left_alpha[17][25] = 1'b1; \
	doodle_left_alpha[17][26] = 1'b1; \
	doodle_left_alpha[17][27] = 1'b1; \
	doodle_left_alpha[17][28] = 1'b1; \
	doodle_left_alpha[17][29] = 1'b1; \
	doodle_left_alpha[17][30] = 1'b1; \
	doodle_left_alpha[17][31] = 1'b0; \
	doodle_left_alpha[17][32] = 1'b0; \
	doodle_left_alpha[17][33] = 1'b0; \
	doodle_left_alpha[17][34] = 1'b0; \
	doodle_left_alpha[17][35] = 1'b0; \
	doodle_left_alpha[17][36] = 1'b0; \
	doodle_left_alpha[17][37] = 1'b0; \
	doodle_left_alpha[17][38] = 1'b0; \
	doodle_left_alpha[17][39] = 1'b0; \
	doodle_left_alpha[17][40] = 1'b0; \
	doodle_left_alpha[17][41] = 1'b0; \
	doodle_left_alpha[17][42] = 1'b0; \
	doodle_left_alpha[17][43] = 1'b0; \
	doodle_left_alpha[17][44] = 1'b0; \
	doodle_left_alpha[17][45] = 1'b0; \
	doodle_left_alpha[17][46] = 1'b0; \
	doodle_left_alpha[17][47] = 1'b0; \
	doodle_left_alpha[17][48] = 1'b0; \
	doodle_left_alpha[17][49] = 1'b0; \
	doodle_left_alpha[17][50] = 1'b0; \
	doodle_left_alpha[17][51] = 1'b0; \
	doodle_left_alpha[17][52] = 1'b0; \
	doodle_left_alpha[17][53] = 1'b0; \
	doodle_left_alpha[17][54] = 1'b0; \
	doodle_left_alpha[17][55] = 1'b0; \
	doodle_left_alpha[17][56] = 1'b0; \
	doodle_left_alpha[17][57] = 1'b1; \
	doodle_left_alpha[17][58] = 1'b1; \
	doodle_left_alpha[17][59] = 1'b1; \
	doodle_left_alpha[17][60] = 1'b1; \
	doodle_left_alpha[17][61] = 1'b1; \
	doodle_left_alpha[17][62] = 1'b1; \
	doodle_left_alpha[17][63] = 1'b1; \
	doodle_left_alpha[17][64] = 1'b1; \
	doodle_left_alpha[17][65] = 1'b1; \
	doodle_left_alpha[17][66] = 1'b1; \
	doodle_left_alpha[17][67] = 1'b1; \
	doodle_left_alpha[17][68] = 1'b1; \
	doodle_left_alpha[17][69] = 1'b1; \
	doodle_left_alpha[17][70] = 1'b1; \
	doodle_left_alpha[17][71] = 1'b1; \
	doodle_left_alpha[17][72] = 1'b1; \
	doodle_left_alpha[17][73] = 1'b1; \
	doodle_left_alpha[17][74] = 1'b1; \
	doodle_left_alpha[17][75] = 1'b1; \
	doodle_left_alpha[17][76] = 1'b1; \
	doodle_left_alpha[17][77] = 1'b1; \
	doodle_left_alpha[17][78] = 1'b1; \
	doodle_left_alpha[17][79] = 1'b1; \
	doodle_left_alpha[18][0] = 1'b1; \
	doodle_left_alpha[18][1] = 1'b1; \
	doodle_left_alpha[18][2] = 1'b1; \
	doodle_left_alpha[18][3] = 1'b1; \
	doodle_left_alpha[18][4] = 1'b1; \
	doodle_left_alpha[18][5] = 1'b1; \
	doodle_left_alpha[18][6] = 1'b1; \
	doodle_left_alpha[18][7] = 1'b1; \
	doodle_left_alpha[18][8] = 1'b1; \
	doodle_left_alpha[18][9] = 1'b1; \
	doodle_left_alpha[18][10] = 1'b1; \
	doodle_left_alpha[18][11] = 1'b1; \
	doodle_left_alpha[18][12] = 1'b1; \
	doodle_left_alpha[18][13] = 1'b1; \
	doodle_left_alpha[18][14] = 1'b1; \
	doodle_left_alpha[18][15] = 1'b1; \
	doodle_left_alpha[18][16] = 1'b1; \
	doodle_left_alpha[18][17] = 1'b1; \
	doodle_left_alpha[18][18] = 1'b1; \
	doodle_left_alpha[18][19] = 1'b1; \
	doodle_left_alpha[18][20] = 1'b1; \
	doodle_left_alpha[18][21] = 1'b1; \
	doodle_left_alpha[18][22] = 1'b1; \
	doodle_left_alpha[18][23] = 1'b1; \
	doodle_left_alpha[18][24] = 1'b1; \
	doodle_left_alpha[18][25] = 1'b1; \
	doodle_left_alpha[18][26] = 1'b1; \
	doodle_left_alpha[18][27] = 1'b1; \
	doodle_left_alpha[18][28] = 1'b1; \
	doodle_left_alpha[18][29] = 1'b1; \
	doodle_left_alpha[18][30] = 1'b1; \
	doodle_left_alpha[18][31] = 1'b0; \
	doodle_left_alpha[18][32] = 1'b0; \
	doodle_left_alpha[18][33] = 1'b0; \
	doodle_left_alpha[18][34] = 1'b0; \
	doodle_left_alpha[18][35] = 1'b0; \
	doodle_left_alpha[18][36] = 1'b0; \
	doodle_left_alpha[18][37] = 1'b0; \
	doodle_left_alpha[18][38] = 1'b0; \
	doodle_left_alpha[18][39] = 1'b0; \
	doodle_left_alpha[18][40] = 1'b0; \
	doodle_left_alpha[18][41] = 1'b0; \
	doodle_left_alpha[18][42] = 1'b0; \
	doodle_left_alpha[18][43] = 1'b0; \
	doodle_left_alpha[18][44] = 1'b0; \
	doodle_left_alpha[18][45] = 1'b0; \
	doodle_left_alpha[18][46] = 1'b0; \
	doodle_left_alpha[18][47] = 1'b0; \
	doodle_left_alpha[18][48] = 1'b0; \
	doodle_left_alpha[18][49] = 1'b0; \
	doodle_left_alpha[18][50] = 1'b0; \
	doodle_left_alpha[18][51] = 1'b0; \
	doodle_left_alpha[18][52] = 1'b0; \
	doodle_left_alpha[18][53] = 1'b0; \
	doodle_left_alpha[18][54] = 1'b0; \
	doodle_left_alpha[18][55] = 1'b0; \
	doodle_left_alpha[18][56] = 1'b0; \
	doodle_left_alpha[18][57] = 1'b1; \
	doodle_left_alpha[18][58] = 1'b1; \
	doodle_left_alpha[18][59] = 1'b1; \
	doodle_left_alpha[18][60] = 1'b1; \
	doodle_left_alpha[18][61] = 1'b1; \
	doodle_left_alpha[18][62] = 1'b1; \
	doodle_left_alpha[18][63] = 1'b1; \
	doodle_left_alpha[18][64] = 1'b1; \
	doodle_left_alpha[18][65] = 1'b1; \
	doodle_left_alpha[18][66] = 1'b1; \
	doodle_left_alpha[18][67] = 1'b1; \
	doodle_left_alpha[18][68] = 1'b1; \
	doodle_left_alpha[18][69] = 1'b1; \
	doodle_left_alpha[18][70] = 1'b1; \
	doodle_left_alpha[18][71] = 1'b1; \
	doodle_left_alpha[18][72] = 1'b1; \
	doodle_left_alpha[18][73] = 1'b1; \
	doodle_left_alpha[18][74] = 1'b1; \
	doodle_left_alpha[18][75] = 1'b1; \
	doodle_left_alpha[18][76] = 1'b1; \
	doodle_left_alpha[18][77] = 1'b1; \
	doodle_left_alpha[18][78] = 1'b1; \
	doodle_left_alpha[18][79] = 1'b1; \
	doodle_left_alpha[19][0] = 1'b1; \
	doodle_left_alpha[19][1] = 1'b1; \
	doodle_left_alpha[19][2] = 1'b1; \
	doodle_left_alpha[19][3] = 1'b1; \
	doodle_left_alpha[19][4] = 1'b1; \
	doodle_left_alpha[19][5] = 1'b1; \
	doodle_left_alpha[19][6] = 1'b1; \
	doodle_left_alpha[19][7] = 1'b1; \
	doodle_left_alpha[19][8] = 1'b1; \
	doodle_left_alpha[19][9] = 1'b1; \
	doodle_left_alpha[19][10] = 1'b1; \
	doodle_left_alpha[19][11] = 1'b1; \
	doodle_left_alpha[19][12] = 1'b1; \
	doodle_left_alpha[19][13] = 1'b1; \
	doodle_left_alpha[19][14] = 1'b1; \
	doodle_left_alpha[19][15] = 1'b1; \
	doodle_left_alpha[19][16] = 1'b1; \
	doodle_left_alpha[19][17] = 1'b1; \
	doodle_left_alpha[19][18] = 1'b1; \
	doodle_left_alpha[19][19] = 1'b1; \
	doodle_left_alpha[19][20] = 1'b1; \
	doodle_left_alpha[19][21] = 1'b1; \
	doodle_left_alpha[19][22] = 1'b1; \
	doodle_left_alpha[19][23] = 1'b1; \
	doodle_left_alpha[19][24] = 1'b1; \
	doodle_left_alpha[19][25] = 1'b1; \
	doodle_left_alpha[19][26] = 1'b1; \
	doodle_left_alpha[19][27] = 1'b1; \
	doodle_left_alpha[19][28] = 1'b1; \
	doodle_left_alpha[19][29] = 1'b1; \
	doodle_left_alpha[19][30] = 1'b1; \
	doodle_left_alpha[19][31] = 1'b0; \
	doodle_left_alpha[19][32] = 1'b0; \
	doodle_left_alpha[19][33] = 1'b0; \
	doodle_left_alpha[19][34] = 1'b0; \
	doodle_left_alpha[19][35] = 1'b0; \
	doodle_left_alpha[19][36] = 1'b0; \
	doodle_left_alpha[19][37] = 1'b0; \
	doodle_left_alpha[19][38] = 1'b0; \
	doodle_left_alpha[19][39] = 1'b0; \
	doodle_left_alpha[19][40] = 1'b0; \
	doodle_left_alpha[19][41] = 1'b0; \
	doodle_left_alpha[19][42] = 1'b0; \
	doodle_left_alpha[19][43] = 1'b0; \
	doodle_left_alpha[19][44] = 1'b0; \
	doodle_left_alpha[19][45] = 1'b0; \
	doodle_left_alpha[19][46] = 1'b0; \
	doodle_left_alpha[19][47] = 1'b0; \
	doodle_left_alpha[19][48] = 1'b0; \
	doodle_left_alpha[19][49] = 1'b0; \
	doodle_left_alpha[19][50] = 1'b0; \
	doodle_left_alpha[19][51] = 1'b0; \
	doodle_left_alpha[19][52] = 1'b0; \
	doodle_left_alpha[19][53] = 1'b0; \
	doodle_left_alpha[19][54] = 1'b0; \
	doodle_left_alpha[19][55] = 1'b0; \
	doodle_left_alpha[19][56] = 1'b0; \
	doodle_left_alpha[19][57] = 1'b1; \
	doodle_left_alpha[19][58] = 1'b1; \
	doodle_left_alpha[19][59] = 1'b1; \
	doodle_left_alpha[19][60] = 1'b1; \
	doodle_left_alpha[19][61] = 1'b1; \
	doodle_left_alpha[19][62] = 1'b1; \
	doodle_left_alpha[19][63] = 1'b1; \
	doodle_left_alpha[19][64] = 1'b1; \
	doodle_left_alpha[19][65] = 1'b1; \
	doodle_left_alpha[19][66] = 1'b1; \
	doodle_left_alpha[19][67] = 1'b1; \
	doodle_left_alpha[19][68] = 1'b1; \
	doodle_left_alpha[19][69] = 1'b1; \
	doodle_left_alpha[19][70] = 1'b1; \
	doodle_left_alpha[19][71] = 1'b1; \
	doodle_left_alpha[19][72] = 1'b1; \
	doodle_left_alpha[19][73] = 1'b1; \
	doodle_left_alpha[19][74] = 1'b1; \
	doodle_left_alpha[19][75] = 1'b1; \
	doodle_left_alpha[19][76] = 1'b1; \
	doodle_left_alpha[19][77] = 1'b1; \
	doodle_left_alpha[19][78] = 1'b1; \
	doodle_left_alpha[19][79] = 1'b1; \
	doodle_left_alpha[20][0] = 1'b1; \
	doodle_left_alpha[20][1] = 1'b1; \
	doodle_left_alpha[20][2] = 1'b1; \
	doodle_left_alpha[20][3] = 1'b1; \
	doodle_left_alpha[20][4] = 1'b1; \
	doodle_left_alpha[20][5] = 1'b1; \
	doodle_left_alpha[20][6] = 1'b1; \
	doodle_left_alpha[20][7] = 1'b1; \
	doodle_left_alpha[20][8] = 1'b1; \
	doodle_left_alpha[20][9] = 1'b1; \
	doodle_left_alpha[20][10] = 1'b1; \
	doodle_left_alpha[20][11] = 1'b1; \
	doodle_left_alpha[20][12] = 1'b1; \
	doodle_left_alpha[20][13] = 1'b1; \
	doodle_left_alpha[20][14] = 1'b1; \
	doodle_left_alpha[20][15] = 1'b1; \
	doodle_left_alpha[20][16] = 1'b1; \
	doodle_left_alpha[20][17] = 1'b1; \
	doodle_left_alpha[20][18] = 1'b1; \
	doodle_left_alpha[20][19] = 1'b1; \
	doodle_left_alpha[20][20] = 1'b1; \
	doodle_left_alpha[20][21] = 1'b1; \
	doodle_left_alpha[20][22] = 1'b1; \
	doodle_left_alpha[20][23] = 1'b1; \
	doodle_left_alpha[20][24] = 1'b1; \
	doodle_left_alpha[20][25] = 1'b1; \
	doodle_left_alpha[20][26] = 1'b1; \
	doodle_left_alpha[20][27] = 1'b0; \
	doodle_left_alpha[20][28] = 1'b0; \
	doodle_left_alpha[20][29] = 1'b0; \
	doodle_left_alpha[20][30] = 1'b0; \
	doodle_left_alpha[20][31] = 1'b0; \
	doodle_left_alpha[20][32] = 1'b0; \
	doodle_left_alpha[20][33] = 1'b0; \
	doodle_left_alpha[20][34] = 1'b0; \
	doodle_left_alpha[20][35] = 1'b0; \
	doodle_left_alpha[20][36] = 1'b0; \
	doodle_left_alpha[20][37] = 1'b0; \
	doodle_left_alpha[20][38] = 1'b0; \
	doodle_left_alpha[20][39] = 1'b0; \
	doodle_left_alpha[20][40] = 1'b0; \
	doodle_left_alpha[20][41] = 1'b0; \
	doodle_left_alpha[20][42] = 1'b0; \
	doodle_left_alpha[20][43] = 1'b0; \
	doodle_left_alpha[20][44] = 1'b0; \
	doodle_left_alpha[20][45] = 1'b0; \
	doodle_left_alpha[20][46] = 1'b0; \
	doodle_left_alpha[20][47] = 1'b0; \
	doodle_left_alpha[20][48] = 1'b0; \
	doodle_left_alpha[20][49] = 1'b0; \
	doodle_left_alpha[20][50] = 1'b0; \
	doodle_left_alpha[20][51] = 1'b0; \
	doodle_left_alpha[20][52] = 1'b0; \
	doodle_left_alpha[20][53] = 1'b0; \
	doodle_left_alpha[20][54] = 1'b0; \
	doodle_left_alpha[20][55] = 1'b0; \
	doodle_left_alpha[20][56] = 1'b0; \
	doodle_left_alpha[20][57] = 1'b0; \
	doodle_left_alpha[20][58] = 1'b0; \
	doodle_left_alpha[20][59] = 1'b0; \
	doodle_left_alpha[20][60] = 1'b0; \
	doodle_left_alpha[20][61] = 1'b1; \
	doodle_left_alpha[20][62] = 1'b1; \
	doodle_left_alpha[20][63] = 1'b1; \
	doodle_left_alpha[20][64] = 1'b1; \
	doodle_left_alpha[20][65] = 1'b1; \
	doodle_left_alpha[20][66] = 1'b1; \
	doodle_left_alpha[20][67] = 1'b1; \
	doodle_left_alpha[20][68] = 1'b1; \
	doodle_left_alpha[20][69] = 1'b1; \
	doodle_left_alpha[20][70] = 1'b1; \
	doodle_left_alpha[20][71] = 1'b1; \
	doodle_left_alpha[20][72] = 1'b1; \
	doodle_left_alpha[20][73] = 1'b1; \
	doodle_left_alpha[20][74] = 1'b1; \
	doodle_left_alpha[20][75] = 1'b1; \
	doodle_left_alpha[20][76] = 1'b1; \
	doodle_left_alpha[20][77] = 1'b1; \
	doodle_left_alpha[20][78] = 1'b1; \
	doodle_left_alpha[20][79] = 1'b1; \
	doodle_left_alpha[21][0] = 1'b1; \
	doodle_left_alpha[21][1] = 1'b1; \
	doodle_left_alpha[21][2] = 1'b1; \
	doodle_left_alpha[21][3] = 1'b1; \
	doodle_left_alpha[21][4] = 1'b1; \
	doodle_left_alpha[21][5] = 1'b1; \
	doodle_left_alpha[21][6] = 1'b1; \
	doodle_left_alpha[21][7] = 1'b1; \
	doodle_left_alpha[21][8] = 1'b1; \
	doodle_left_alpha[21][9] = 1'b1; \
	doodle_left_alpha[21][10] = 1'b1; \
	doodle_left_alpha[21][11] = 1'b1; \
	doodle_left_alpha[21][12] = 1'b1; \
	doodle_left_alpha[21][13] = 1'b1; \
	doodle_left_alpha[21][14] = 1'b1; \
	doodle_left_alpha[21][15] = 1'b1; \
	doodle_left_alpha[21][16] = 1'b1; \
	doodle_left_alpha[21][17] = 1'b1; \
	doodle_left_alpha[21][18] = 1'b1; \
	doodle_left_alpha[21][19] = 1'b1; \
	doodle_left_alpha[21][20] = 1'b1; \
	doodle_left_alpha[21][21] = 1'b1; \
	doodle_left_alpha[21][22] = 1'b1; \
	doodle_left_alpha[21][23] = 1'b1; \
	doodle_left_alpha[21][24] = 1'b1; \
	doodle_left_alpha[21][25] = 1'b1; \
	doodle_left_alpha[21][26] = 1'b1; \
	doodle_left_alpha[21][27] = 1'b0; \
	doodle_left_alpha[21][28] = 1'b0; \
	doodle_left_alpha[21][29] = 1'b0; \
	doodle_left_alpha[21][30] = 1'b0; \
	doodle_left_alpha[21][31] = 1'b0; \
	doodle_left_alpha[21][32] = 1'b0; \
	doodle_left_alpha[21][33] = 1'b0; \
	doodle_left_alpha[21][34] = 1'b0; \
	doodle_left_alpha[21][35] = 1'b0; \
	doodle_left_alpha[21][36] = 1'b0; \
	doodle_left_alpha[21][37] = 1'b0; \
	doodle_left_alpha[21][38] = 1'b0; \
	doodle_left_alpha[21][39] = 1'b0; \
	doodle_left_alpha[21][40] = 1'b0; \
	doodle_left_alpha[21][41] = 1'b0; \
	doodle_left_alpha[21][42] = 1'b0; \
	doodle_left_alpha[21][43] = 1'b0; \
	doodle_left_alpha[21][44] = 1'b0; \
	doodle_left_alpha[21][45] = 1'b0; \
	doodle_left_alpha[21][46] = 1'b0; \
	doodle_left_alpha[21][47] = 1'b0; \
	doodle_left_alpha[21][48] = 1'b0; \
	doodle_left_alpha[21][49] = 1'b0; \
	doodle_left_alpha[21][50] = 1'b0; \
	doodle_left_alpha[21][51] = 1'b0; \
	doodle_left_alpha[21][52] = 1'b0; \
	doodle_left_alpha[21][53] = 1'b0; \
	doodle_left_alpha[21][54] = 1'b0; \
	doodle_left_alpha[21][55] = 1'b0; \
	doodle_left_alpha[21][56] = 1'b0; \
	doodle_left_alpha[21][57] = 1'b0; \
	doodle_left_alpha[21][58] = 1'b0; \
	doodle_left_alpha[21][59] = 1'b0; \
	doodle_left_alpha[21][60] = 1'b0; \
	doodle_left_alpha[21][61] = 1'b1; \
	doodle_left_alpha[21][62] = 1'b1; \
	doodle_left_alpha[21][63] = 1'b1; \
	doodle_left_alpha[21][64] = 1'b1; \
	doodle_left_alpha[21][65] = 1'b1; \
	doodle_left_alpha[21][66] = 1'b1; \
	doodle_left_alpha[21][67] = 1'b1; \
	doodle_left_alpha[21][68] = 1'b1; \
	doodle_left_alpha[21][69] = 1'b1; \
	doodle_left_alpha[21][70] = 1'b1; \
	doodle_left_alpha[21][71] = 1'b1; \
	doodle_left_alpha[21][72] = 1'b1; \
	doodle_left_alpha[21][73] = 1'b1; \
	doodle_left_alpha[21][74] = 1'b1; \
	doodle_left_alpha[21][75] = 1'b1; \
	doodle_left_alpha[21][76] = 1'b1; \
	doodle_left_alpha[21][77] = 1'b1; \
	doodle_left_alpha[21][78] = 1'b1; \
	doodle_left_alpha[21][79] = 1'b1; \
	doodle_left_alpha[22][0] = 1'b1; \
	doodle_left_alpha[22][1] = 1'b1; \
	doodle_left_alpha[22][2] = 1'b1; \
	doodle_left_alpha[22][3] = 1'b1; \
	doodle_left_alpha[22][4] = 1'b1; \
	doodle_left_alpha[22][5] = 1'b1; \
	doodle_left_alpha[22][6] = 1'b1; \
	doodle_left_alpha[22][7] = 1'b1; \
	doodle_left_alpha[22][8] = 1'b1; \
	doodle_left_alpha[22][9] = 1'b1; \
	doodle_left_alpha[22][10] = 1'b1; \
	doodle_left_alpha[22][11] = 1'b1; \
	doodle_left_alpha[22][12] = 1'b1; \
	doodle_left_alpha[22][13] = 1'b1; \
	doodle_left_alpha[22][14] = 1'b1; \
	doodle_left_alpha[22][15] = 1'b1; \
	doodle_left_alpha[22][16] = 1'b1; \
	doodle_left_alpha[22][17] = 1'b1; \
	doodle_left_alpha[22][18] = 1'b1; \
	doodle_left_alpha[22][19] = 1'b1; \
	doodle_left_alpha[22][20] = 1'b1; \
	doodle_left_alpha[22][21] = 1'b1; \
	doodle_left_alpha[22][22] = 1'b1; \
	doodle_left_alpha[22][23] = 1'b1; \
	doodle_left_alpha[22][24] = 1'b1; \
	doodle_left_alpha[22][25] = 1'b1; \
	doodle_left_alpha[22][26] = 1'b1; \
	doodle_left_alpha[22][27] = 1'b0; \
	doodle_left_alpha[22][28] = 1'b0; \
	doodle_left_alpha[22][29] = 1'b0; \
	doodle_left_alpha[22][30] = 1'b0; \
	doodle_left_alpha[22][31] = 1'b0; \
	doodle_left_alpha[22][32] = 1'b0; \
	doodle_left_alpha[22][33] = 1'b0; \
	doodle_left_alpha[22][34] = 1'b0; \
	doodle_left_alpha[22][35] = 1'b0; \
	doodle_left_alpha[22][36] = 1'b0; \
	doodle_left_alpha[22][37] = 1'b0; \
	doodle_left_alpha[22][38] = 1'b0; \
	doodle_left_alpha[22][39] = 1'b0; \
	doodle_left_alpha[22][40] = 1'b0; \
	doodle_left_alpha[22][41] = 1'b0; \
	doodle_left_alpha[22][42] = 1'b0; \
	doodle_left_alpha[22][43] = 1'b0; \
	doodle_left_alpha[22][44] = 1'b0; \
	doodle_left_alpha[22][45] = 1'b0; \
	doodle_left_alpha[22][46] = 1'b0; \
	doodle_left_alpha[22][47] = 1'b0; \
	doodle_left_alpha[22][48] = 1'b0; \
	doodle_left_alpha[22][49] = 1'b0; \
	doodle_left_alpha[22][50] = 1'b0; \
	doodle_left_alpha[22][51] = 1'b0; \
	doodle_left_alpha[22][52] = 1'b0; \
	doodle_left_alpha[22][53] = 1'b0; \
	doodle_left_alpha[22][54] = 1'b0; \
	doodle_left_alpha[22][55] = 1'b0; \
	doodle_left_alpha[22][56] = 1'b0; \
	doodle_left_alpha[22][57] = 1'b0; \
	doodle_left_alpha[22][58] = 1'b0; \
	doodle_left_alpha[22][59] = 1'b0; \
	doodle_left_alpha[22][60] = 1'b0; \
	doodle_left_alpha[22][61] = 1'b1; \
	doodle_left_alpha[22][62] = 1'b1; \
	doodle_left_alpha[22][63] = 1'b1; \
	doodle_left_alpha[22][64] = 1'b1; \
	doodle_left_alpha[22][65] = 1'b1; \
	doodle_left_alpha[22][66] = 1'b1; \
	doodle_left_alpha[22][67] = 1'b1; \
	doodle_left_alpha[22][68] = 1'b1; \
	doodle_left_alpha[22][69] = 1'b1; \
	doodle_left_alpha[22][70] = 1'b1; \
	doodle_left_alpha[22][71] = 1'b1; \
	doodle_left_alpha[22][72] = 1'b1; \
	doodle_left_alpha[22][73] = 1'b1; \
	doodle_left_alpha[22][74] = 1'b1; \
	doodle_left_alpha[22][75] = 1'b1; \
	doodle_left_alpha[22][76] = 1'b1; \
	doodle_left_alpha[22][77] = 1'b1; \
	doodle_left_alpha[22][78] = 1'b1; \
	doodle_left_alpha[22][79] = 1'b1; \
	doodle_left_alpha[23][0] = 1'b1; \
	doodle_left_alpha[23][1] = 1'b1; \
	doodle_left_alpha[23][2] = 1'b1; \
	doodle_left_alpha[23][3] = 1'b1; \
	doodle_left_alpha[23][4] = 1'b1; \
	doodle_left_alpha[23][5] = 1'b1; \
	doodle_left_alpha[23][6] = 1'b1; \
	doodle_left_alpha[23][7] = 1'b1; \
	doodle_left_alpha[23][8] = 1'b1; \
	doodle_left_alpha[23][9] = 1'b1; \
	doodle_left_alpha[23][10] = 1'b1; \
	doodle_left_alpha[23][11] = 1'b1; \
	doodle_left_alpha[23][12] = 1'b1; \
	doodle_left_alpha[23][13] = 1'b1; \
	doodle_left_alpha[23][14] = 1'b1; \
	doodle_left_alpha[23][15] = 1'b1; \
	doodle_left_alpha[23][16] = 1'b1; \
	doodle_left_alpha[23][17] = 1'b1; \
	doodle_left_alpha[23][18] = 1'b1; \
	doodle_left_alpha[23][19] = 1'b1; \
	doodle_left_alpha[23][20] = 1'b1; \
	doodle_left_alpha[23][21] = 1'b1; \
	doodle_left_alpha[23][22] = 1'b1; \
	doodle_left_alpha[23][23] = 1'b1; \
	doodle_left_alpha[23][24] = 1'b1; \
	doodle_left_alpha[23][25] = 1'b1; \
	doodle_left_alpha[23][26] = 1'b1; \
	doodle_left_alpha[23][27] = 1'b0; \
	doodle_left_alpha[23][28] = 1'b0; \
	doodle_left_alpha[23][29] = 1'b0; \
	doodle_left_alpha[23][30] = 1'b0; \
	doodle_left_alpha[23][31] = 1'b0; \
	doodle_left_alpha[23][32] = 1'b0; \
	doodle_left_alpha[23][33] = 1'b0; \
	doodle_left_alpha[23][34] = 1'b0; \
	doodle_left_alpha[23][35] = 1'b0; \
	doodle_left_alpha[23][36] = 1'b0; \
	doodle_left_alpha[23][37] = 1'b0; \
	doodle_left_alpha[23][38] = 1'b0; \
	doodle_left_alpha[23][39] = 1'b0; \
	doodle_left_alpha[23][40] = 1'b0; \
	doodle_left_alpha[23][41] = 1'b0; \
	doodle_left_alpha[23][42] = 1'b0; \
	doodle_left_alpha[23][43] = 1'b0; \
	doodle_left_alpha[23][44] = 1'b0; \
	doodle_left_alpha[23][45] = 1'b0; \
	doodle_left_alpha[23][46] = 1'b0; \
	doodle_left_alpha[23][47] = 1'b0; \
	doodle_left_alpha[23][48] = 1'b0; \
	doodle_left_alpha[23][49] = 1'b0; \
	doodle_left_alpha[23][50] = 1'b0; \
	doodle_left_alpha[23][51] = 1'b0; \
	doodle_left_alpha[23][52] = 1'b0; \
	doodle_left_alpha[23][53] = 1'b0; \
	doodle_left_alpha[23][54] = 1'b0; \
	doodle_left_alpha[23][55] = 1'b0; \
	doodle_left_alpha[23][56] = 1'b0; \
	doodle_left_alpha[23][57] = 1'b0; \
	doodle_left_alpha[23][58] = 1'b0; \
	doodle_left_alpha[23][59] = 1'b0; \
	doodle_left_alpha[23][60] = 1'b0; \
	doodle_left_alpha[23][61] = 1'b1; \
	doodle_left_alpha[23][62] = 1'b1; \
	doodle_left_alpha[23][63] = 1'b1; \
	doodle_left_alpha[23][64] = 1'b1; \
	doodle_left_alpha[23][65] = 1'b1; \
	doodle_left_alpha[23][66] = 1'b1; \
	doodle_left_alpha[23][67] = 1'b1; \
	doodle_left_alpha[23][68] = 1'b1; \
	doodle_left_alpha[23][69] = 1'b1; \
	doodle_left_alpha[23][70] = 1'b1; \
	doodle_left_alpha[23][71] = 1'b1; \
	doodle_left_alpha[23][72] = 1'b1; \
	doodle_left_alpha[23][73] = 1'b1; \
	doodle_left_alpha[23][74] = 1'b1; \
	doodle_left_alpha[23][75] = 1'b1; \
	doodle_left_alpha[23][76] = 1'b1; \
	doodle_left_alpha[23][77] = 1'b1; \
	doodle_left_alpha[23][78] = 1'b1; \
	doodle_left_alpha[23][79] = 1'b1; \
	doodle_left_alpha[24][0] = 1'b1; \
	doodle_left_alpha[24][1] = 1'b1; \
	doodle_left_alpha[24][2] = 1'b1; \
	doodle_left_alpha[24][3] = 1'b1; \
	doodle_left_alpha[24][4] = 1'b1; \
	doodle_left_alpha[24][5] = 1'b1; \
	doodle_left_alpha[24][6] = 1'b1; \
	doodle_left_alpha[24][7] = 1'b1; \
	doodle_left_alpha[24][8] = 1'b1; \
	doodle_left_alpha[24][9] = 1'b1; \
	doodle_left_alpha[24][10] = 1'b1; \
	doodle_left_alpha[24][11] = 1'b1; \
	doodle_left_alpha[24][12] = 1'b1; \
	doodle_left_alpha[24][13] = 1'b1; \
	doodle_left_alpha[24][14] = 1'b1; \
	doodle_left_alpha[24][15] = 1'b1; \
	doodle_left_alpha[24][16] = 1'b1; \
	doodle_left_alpha[24][17] = 1'b1; \
	doodle_left_alpha[24][18] = 1'b1; \
	doodle_left_alpha[24][19] = 1'b1; \
	doodle_left_alpha[24][20] = 1'b1; \
	doodle_left_alpha[24][21] = 1'b1; \
	doodle_left_alpha[24][22] = 1'b1; \
	doodle_left_alpha[24][23] = 1'b0; \
	doodle_left_alpha[24][24] = 1'b0; \
	doodle_left_alpha[24][25] = 1'b0; \
	doodle_left_alpha[24][26] = 1'b0; \
	doodle_left_alpha[24][27] = 1'b0; \
	doodle_left_alpha[24][28] = 1'b0; \
	doodle_left_alpha[24][29] = 1'b0; \
	doodle_left_alpha[24][30] = 1'b0; \
	doodle_left_alpha[24][31] = 1'b0; \
	doodle_left_alpha[24][32] = 1'b0; \
	doodle_left_alpha[24][33] = 1'b0; \
	doodle_left_alpha[24][34] = 1'b0; \
	doodle_left_alpha[24][35] = 1'b0; \
	doodle_left_alpha[24][36] = 1'b0; \
	doodle_left_alpha[24][37] = 1'b0; \
	doodle_left_alpha[24][38] = 1'b0; \
	doodle_left_alpha[24][39] = 1'b0; \
	doodle_left_alpha[24][40] = 1'b0; \
	doodle_left_alpha[24][41] = 1'b0; \
	doodle_left_alpha[24][42] = 1'b0; \
	doodle_left_alpha[24][43] = 1'b0; \
	doodle_left_alpha[24][44] = 1'b0; \
	doodle_left_alpha[24][45] = 1'b0; \
	doodle_left_alpha[24][46] = 1'b0; \
	doodle_left_alpha[24][47] = 1'b0; \
	doodle_left_alpha[24][48] = 1'b0; \
	doodle_left_alpha[24][49] = 1'b0; \
	doodle_left_alpha[24][50] = 1'b0; \
	doodle_left_alpha[24][51] = 1'b0; \
	doodle_left_alpha[24][52] = 1'b0; \
	doodle_left_alpha[24][53] = 1'b0; \
	doodle_left_alpha[24][54] = 1'b0; \
	doodle_left_alpha[24][55] = 1'b0; \
	doodle_left_alpha[24][56] = 1'b0; \
	doodle_left_alpha[24][57] = 1'b0; \
	doodle_left_alpha[24][58] = 1'b0; \
	doodle_left_alpha[24][59] = 1'b0; \
	doodle_left_alpha[24][60] = 1'b0; \
	doodle_left_alpha[24][61] = 1'b0; \
	doodle_left_alpha[24][62] = 1'b0; \
	doodle_left_alpha[24][63] = 1'b0; \
	doodle_left_alpha[24][64] = 1'b0; \
	doodle_left_alpha[24][65] = 1'b1; \
	doodle_left_alpha[24][66] = 1'b1; \
	doodle_left_alpha[24][67] = 1'b1; \
	doodle_left_alpha[24][68] = 1'b1; \
	doodle_left_alpha[24][69] = 1'b1; \
	doodle_left_alpha[24][70] = 1'b1; \
	doodle_left_alpha[24][71] = 1'b1; \
	doodle_left_alpha[24][72] = 1'b1; \
	doodle_left_alpha[24][73] = 1'b1; \
	doodle_left_alpha[24][74] = 1'b1; \
	doodle_left_alpha[24][75] = 1'b1; \
	doodle_left_alpha[24][76] = 1'b1; \
	doodle_left_alpha[24][77] = 1'b1; \
	doodle_left_alpha[24][78] = 1'b1; \
	doodle_left_alpha[24][79] = 1'b1; \
	doodle_left_alpha[25][0] = 1'b1; \
	doodle_left_alpha[25][1] = 1'b1; \
	doodle_left_alpha[25][2] = 1'b1; \
	doodle_left_alpha[25][3] = 1'b1; \
	doodle_left_alpha[25][4] = 1'b1; \
	doodle_left_alpha[25][5] = 1'b1; \
	doodle_left_alpha[25][6] = 1'b1; \
	doodle_left_alpha[25][7] = 1'b1; \
	doodle_left_alpha[25][8] = 1'b1; \
	doodle_left_alpha[25][9] = 1'b1; \
	doodle_left_alpha[25][10] = 1'b1; \
	doodle_left_alpha[25][11] = 1'b1; \
	doodle_left_alpha[25][12] = 1'b1; \
	doodle_left_alpha[25][13] = 1'b1; \
	doodle_left_alpha[25][14] = 1'b1; \
	doodle_left_alpha[25][15] = 1'b1; \
	doodle_left_alpha[25][16] = 1'b1; \
	doodle_left_alpha[25][17] = 1'b1; \
	doodle_left_alpha[25][18] = 1'b1; \
	doodle_left_alpha[25][19] = 1'b1; \
	doodle_left_alpha[25][20] = 1'b1; \
	doodle_left_alpha[25][21] = 1'b1; \
	doodle_left_alpha[25][22] = 1'b1; \
	doodle_left_alpha[25][23] = 1'b0; \
	doodle_left_alpha[25][24] = 1'b0; \
	doodle_left_alpha[25][25] = 1'b0; \
	doodle_left_alpha[25][26] = 1'b0; \
	doodle_left_alpha[25][27] = 1'b0; \
	doodle_left_alpha[25][28] = 1'b0; \
	doodle_left_alpha[25][29] = 1'b0; \
	doodle_left_alpha[25][30] = 1'b0; \
	doodle_left_alpha[25][31] = 1'b0; \
	doodle_left_alpha[25][32] = 1'b0; \
	doodle_left_alpha[25][33] = 1'b0; \
	doodle_left_alpha[25][34] = 1'b0; \
	doodle_left_alpha[25][35] = 1'b0; \
	doodle_left_alpha[25][36] = 1'b0; \
	doodle_left_alpha[25][37] = 1'b0; \
	doodle_left_alpha[25][38] = 1'b0; \
	doodle_left_alpha[25][39] = 1'b0; \
	doodle_left_alpha[25][40] = 1'b0; \
	doodle_left_alpha[25][41] = 1'b0; \
	doodle_left_alpha[25][42] = 1'b0; \
	doodle_left_alpha[25][43] = 1'b0; \
	doodle_left_alpha[25][44] = 1'b0; \
	doodle_left_alpha[25][45] = 1'b0; \
	doodle_left_alpha[25][46] = 1'b0; \
	doodle_left_alpha[25][47] = 1'b0; \
	doodle_left_alpha[25][48] = 1'b0; \
	doodle_left_alpha[25][49] = 1'b0; \
	doodle_left_alpha[25][50] = 1'b0; \
	doodle_left_alpha[25][51] = 1'b0; \
	doodle_left_alpha[25][52] = 1'b0; \
	doodle_left_alpha[25][53] = 1'b0; \
	doodle_left_alpha[25][54] = 1'b0; \
	doodle_left_alpha[25][55] = 1'b0; \
	doodle_left_alpha[25][56] = 1'b0; \
	doodle_left_alpha[25][57] = 1'b0; \
	doodle_left_alpha[25][58] = 1'b0; \
	doodle_left_alpha[25][59] = 1'b0; \
	doodle_left_alpha[25][60] = 1'b0; \
	doodle_left_alpha[25][61] = 1'b0; \
	doodle_left_alpha[25][62] = 1'b0; \
	doodle_left_alpha[25][63] = 1'b0; \
	doodle_left_alpha[25][64] = 1'b0; \
	doodle_left_alpha[25][65] = 1'b1; \
	doodle_left_alpha[25][66] = 1'b1; \
	doodle_left_alpha[25][67] = 1'b1; \
	doodle_left_alpha[25][68] = 1'b1; \
	doodle_left_alpha[25][69] = 1'b1; \
	doodle_left_alpha[25][70] = 1'b1; \
	doodle_left_alpha[25][71] = 1'b1; \
	doodle_left_alpha[25][72] = 1'b1; \
	doodle_left_alpha[25][73] = 1'b1; \
	doodle_left_alpha[25][74] = 1'b1; \
	doodle_left_alpha[25][75] = 1'b1; \
	doodle_left_alpha[25][76] = 1'b1; \
	doodle_left_alpha[25][77] = 1'b1; \
	doodle_left_alpha[25][78] = 1'b1; \
	doodle_left_alpha[25][79] = 1'b1; \
	doodle_left_alpha[26][0] = 1'b1; \
	doodle_left_alpha[26][1] = 1'b1; \
	doodle_left_alpha[26][2] = 1'b1; \
	doodle_left_alpha[26][3] = 1'b1; \
	doodle_left_alpha[26][4] = 1'b1; \
	doodle_left_alpha[26][5] = 1'b1; \
	doodle_left_alpha[26][6] = 1'b1; \
	doodle_left_alpha[26][7] = 1'b1; \
	doodle_left_alpha[26][8] = 1'b1; \
	doodle_left_alpha[26][9] = 1'b1; \
	doodle_left_alpha[26][10] = 1'b1; \
	doodle_left_alpha[26][11] = 1'b1; \
	doodle_left_alpha[26][12] = 1'b1; \
	doodle_left_alpha[26][13] = 1'b1; \
	doodle_left_alpha[26][14] = 1'b1; \
	doodle_left_alpha[26][15] = 1'b1; \
	doodle_left_alpha[26][16] = 1'b1; \
	doodle_left_alpha[26][17] = 1'b1; \
	doodle_left_alpha[26][18] = 1'b1; \
	doodle_left_alpha[26][19] = 1'b1; \
	doodle_left_alpha[26][20] = 1'b1; \
	doodle_left_alpha[26][21] = 1'b1; \
	doodle_left_alpha[26][22] = 1'b1; \
	doodle_left_alpha[26][23] = 1'b0; \
	doodle_left_alpha[26][24] = 1'b0; \
	doodle_left_alpha[26][25] = 1'b0; \
	doodle_left_alpha[26][26] = 1'b0; \
	doodle_left_alpha[26][27] = 1'b0; \
	doodle_left_alpha[26][28] = 1'b0; \
	doodle_left_alpha[26][29] = 1'b0; \
	doodle_left_alpha[26][30] = 1'b0; \
	doodle_left_alpha[26][31] = 1'b0; \
	doodle_left_alpha[26][32] = 1'b0; \
	doodle_left_alpha[26][33] = 1'b0; \
	doodle_left_alpha[26][34] = 1'b0; \
	doodle_left_alpha[26][35] = 1'b0; \
	doodle_left_alpha[26][36] = 1'b0; \
	doodle_left_alpha[26][37] = 1'b0; \
	doodle_left_alpha[26][38] = 1'b0; \
	doodle_left_alpha[26][39] = 1'b0; \
	doodle_left_alpha[26][40] = 1'b0; \
	doodle_left_alpha[26][41] = 1'b0; \
	doodle_left_alpha[26][42] = 1'b0; \
	doodle_left_alpha[26][43] = 1'b0; \
	doodle_left_alpha[26][44] = 1'b0; \
	doodle_left_alpha[26][45] = 1'b0; \
	doodle_left_alpha[26][46] = 1'b0; \
	doodle_left_alpha[26][47] = 1'b0; \
	doodle_left_alpha[26][48] = 1'b0; \
	doodle_left_alpha[26][49] = 1'b0; \
	doodle_left_alpha[26][50] = 1'b0; \
	doodle_left_alpha[26][51] = 1'b0; \
	doodle_left_alpha[26][52] = 1'b0; \
	doodle_left_alpha[26][53] = 1'b0; \
	doodle_left_alpha[26][54] = 1'b0; \
	doodle_left_alpha[26][55] = 1'b0; \
	doodle_left_alpha[26][56] = 1'b0; \
	doodle_left_alpha[26][57] = 1'b0; \
	doodle_left_alpha[26][58] = 1'b0; \
	doodle_left_alpha[26][59] = 1'b0; \
	doodle_left_alpha[26][60] = 1'b0; \
	doodle_left_alpha[26][61] = 1'b0; \
	doodle_left_alpha[26][62] = 1'b0; \
	doodle_left_alpha[26][63] = 1'b0; \
	doodle_left_alpha[26][64] = 1'b0; \
	doodle_left_alpha[26][65] = 1'b1; \
	doodle_left_alpha[26][66] = 1'b1; \
	doodle_left_alpha[26][67] = 1'b1; \
	doodle_left_alpha[26][68] = 1'b1; \
	doodle_left_alpha[26][69] = 1'b1; \
	doodle_left_alpha[26][70] = 1'b1; \
	doodle_left_alpha[26][71] = 1'b1; \
	doodle_left_alpha[26][72] = 1'b1; \
	doodle_left_alpha[26][73] = 1'b1; \
	doodle_left_alpha[26][74] = 1'b1; \
	doodle_left_alpha[26][75] = 1'b1; \
	doodle_left_alpha[26][76] = 1'b1; \
	doodle_left_alpha[26][77] = 1'b1; \
	doodle_left_alpha[26][78] = 1'b1; \
	doodle_left_alpha[26][79] = 1'b1; \
	doodle_left_alpha[27][0] = 1'b1; \
	doodle_left_alpha[27][1] = 1'b1; \
	doodle_left_alpha[27][2] = 1'b1; \
	doodle_left_alpha[27][3] = 1'b1; \
	doodle_left_alpha[27][4] = 1'b1; \
	doodle_left_alpha[27][5] = 1'b1; \
	doodle_left_alpha[27][6] = 1'b1; \
	doodle_left_alpha[27][7] = 1'b1; \
	doodle_left_alpha[27][8] = 1'b1; \
	doodle_left_alpha[27][9] = 1'b1; \
	doodle_left_alpha[27][10] = 1'b1; \
	doodle_left_alpha[27][11] = 1'b1; \
	doodle_left_alpha[27][12] = 1'b1; \
	doodle_left_alpha[27][13] = 1'b1; \
	doodle_left_alpha[27][14] = 1'b1; \
	doodle_left_alpha[27][15] = 1'b1; \
	doodle_left_alpha[27][16] = 1'b1; \
	doodle_left_alpha[27][17] = 1'b1; \
	doodle_left_alpha[27][18] = 1'b1; \
	doodle_left_alpha[27][19] = 1'b1; \
	doodle_left_alpha[27][20] = 1'b1; \
	doodle_left_alpha[27][21] = 1'b1; \
	doodle_left_alpha[27][22] = 1'b1; \
	doodle_left_alpha[27][23] = 1'b0; \
	doodle_left_alpha[27][24] = 1'b0; \
	doodle_left_alpha[27][25] = 1'b0; \
	doodle_left_alpha[27][26] = 1'b0; \
	doodle_left_alpha[27][27] = 1'b0; \
	doodle_left_alpha[27][28] = 1'b0; \
	doodle_left_alpha[27][29] = 1'b0; \
	doodle_left_alpha[27][30] = 1'b0; \
	doodle_left_alpha[27][31] = 1'b0; \
	doodle_left_alpha[27][32] = 1'b0; \
	doodle_left_alpha[27][33] = 1'b0; \
	doodle_left_alpha[27][34] = 1'b0; \
	doodle_left_alpha[27][35] = 1'b0; \
	doodle_left_alpha[27][36] = 1'b0; \
	doodle_left_alpha[27][37] = 1'b0; \
	doodle_left_alpha[27][38] = 1'b0; \
	doodle_left_alpha[27][39] = 1'b0; \
	doodle_left_alpha[27][40] = 1'b0; \
	doodle_left_alpha[27][41] = 1'b0; \
	doodle_left_alpha[27][42] = 1'b0; \
	doodle_left_alpha[27][43] = 1'b0; \
	doodle_left_alpha[27][44] = 1'b0; \
	doodle_left_alpha[27][45] = 1'b0; \
	doodle_left_alpha[27][46] = 1'b0; \
	doodle_left_alpha[27][47] = 1'b0; \
	doodle_left_alpha[27][48] = 1'b0; \
	doodle_left_alpha[27][49] = 1'b0; \
	doodle_left_alpha[27][50] = 1'b0; \
	doodle_left_alpha[27][51] = 1'b0; \
	doodle_left_alpha[27][52] = 1'b0; \
	doodle_left_alpha[27][53] = 1'b0; \
	doodle_left_alpha[27][54] = 1'b0; \
	doodle_left_alpha[27][55] = 1'b0; \
	doodle_left_alpha[27][56] = 1'b0; \
	doodle_left_alpha[27][57] = 1'b0; \
	doodle_left_alpha[27][58] = 1'b0; \
	doodle_left_alpha[27][59] = 1'b0; \
	doodle_left_alpha[27][60] = 1'b0; \
	doodle_left_alpha[27][61] = 1'b0; \
	doodle_left_alpha[27][62] = 1'b0; \
	doodle_left_alpha[27][63] = 1'b0; \
	doodle_left_alpha[27][64] = 1'b0; \
	doodle_left_alpha[27][65] = 1'b1; \
	doodle_left_alpha[27][66] = 1'b1; \
	doodle_left_alpha[27][67] = 1'b1; \
	doodle_left_alpha[27][68] = 1'b1; \
	doodle_left_alpha[27][69] = 1'b1; \
	doodle_left_alpha[27][70] = 1'b1; \
	doodle_left_alpha[27][71] = 1'b1; \
	doodle_left_alpha[27][72] = 1'b1; \
	doodle_left_alpha[27][73] = 1'b1; \
	doodle_left_alpha[27][74] = 1'b1; \
	doodle_left_alpha[27][75] = 1'b1; \
	doodle_left_alpha[27][76] = 1'b1; \
	doodle_left_alpha[27][77] = 1'b1; \
	doodle_left_alpha[27][78] = 1'b1; \
	doodle_left_alpha[27][79] = 1'b1; \
	doodle_left_alpha[28][0] = 1'b1; \
	doodle_left_alpha[28][1] = 1'b1; \
	doodle_left_alpha[28][2] = 1'b1; \
	doodle_left_alpha[28][3] = 1'b1; \
	doodle_left_alpha[28][4] = 1'b1; \
	doodle_left_alpha[28][5] = 1'b1; \
	doodle_left_alpha[28][6] = 1'b1; \
	doodle_left_alpha[28][7] = 1'b1; \
	doodle_left_alpha[28][8] = 1'b1; \
	doodle_left_alpha[28][9] = 1'b1; \
	doodle_left_alpha[28][10] = 1'b1; \
	doodle_left_alpha[28][11] = 1'b1; \
	doodle_left_alpha[28][12] = 1'b1; \
	doodle_left_alpha[28][13] = 1'b1; \
	doodle_left_alpha[28][14] = 1'b1; \
	doodle_left_alpha[28][15] = 1'b1; \
	doodle_left_alpha[28][16] = 1'b1; \
	doodle_left_alpha[28][17] = 1'b1; \
	doodle_left_alpha[28][18] = 1'b1; \
	doodle_left_alpha[28][19] = 1'b1; \
	doodle_left_alpha[28][20] = 1'b1; \
	doodle_left_alpha[28][21] = 1'b1; \
	doodle_left_alpha[28][22] = 1'b1; \
	doodle_left_alpha[28][23] = 1'b0; \
	doodle_left_alpha[28][24] = 1'b0; \
	doodle_left_alpha[28][25] = 1'b0; \
	doodle_left_alpha[28][26] = 1'b0; \
	doodle_left_alpha[28][27] = 1'b0; \
	doodle_left_alpha[28][28] = 1'b0; \
	doodle_left_alpha[28][29] = 1'b0; \
	doodle_left_alpha[28][30] = 1'b0; \
	doodle_left_alpha[28][31] = 1'b0; \
	doodle_left_alpha[28][32] = 1'b0; \
	doodle_left_alpha[28][33] = 1'b0; \
	doodle_left_alpha[28][34] = 1'b0; \
	doodle_left_alpha[28][35] = 1'b0; \
	doodle_left_alpha[28][36] = 1'b0; \
	doodle_left_alpha[28][37] = 1'b0; \
	doodle_left_alpha[28][38] = 1'b0; \
	doodle_left_alpha[28][39] = 1'b0; \
	doodle_left_alpha[28][40] = 1'b0; \
	doodle_left_alpha[28][41] = 1'b0; \
	doodle_left_alpha[28][42] = 1'b0; \
	doodle_left_alpha[28][43] = 1'b0; \
	doodle_left_alpha[28][44] = 1'b0; \
	doodle_left_alpha[28][45] = 1'b0; \
	doodle_left_alpha[28][46] = 1'b0; \
	doodle_left_alpha[28][47] = 1'b0; \
	doodle_left_alpha[28][48] = 1'b0; \
	doodle_left_alpha[28][49] = 1'b0; \
	doodle_left_alpha[28][50] = 1'b0; \
	doodle_left_alpha[28][51] = 1'b0; \
	doodle_left_alpha[28][52] = 1'b0; \
	doodle_left_alpha[28][53] = 1'b0; \
	doodle_left_alpha[28][54] = 1'b0; \
	doodle_left_alpha[28][55] = 1'b0; \
	doodle_left_alpha[28][56] = 1'b0; \
	doodle_left_alpha[28][57] = 1'b0; \
	doodle_left_alpha[28][58] = 1'b0; \
	doodle_left_alpha[28][59] = 1'b0; \
	doodle_left_alpha[28][60] = 1'b0; \
	doodle_left_alpha[28][61] = 1'b0; \
	doodle_left_alpha[28][62] = 1'b0; \
	doodle_left_alpha[28][63] = 1'b0; \
	doodle_left_alpha[28][64] = 1'b0; \
	doodle_left_alpha[28][65] = 1'b1; \
	doodle_left_alpha[28][66] = 1'b1; \
	doodle_left_alpha[28][67] = 1'b1; \
	doodle_left_alpha[28][68] = 1'b1; \
	doodle_left_alpha[28][69] = 1'b1; \
	doodle_left_alpha[28][70] = 1'b1; \
	doodle_left_alpha[28][71] = 1'b1; \
	doodle_left_alpha[28][72] = 1'b1; \
	doodle_left_alpha[28][73] = 1'b1; \
	doodle_left_alpha[28][74] = 1'b1; \
	doodle_left_alpha[28][75] = 1'b1; \
	doodle_left_alpha[28][76] = 1'b1; \
	doodle_left_alpha[28][77] = 1'b1; \
	doodle_left_alpha[28][78] = 1'b1; \
	doodle_left_alpha[28][79] = 1'b1; \
	doodle_left_alpha[29][0] = 1'b1; \
	doodle_left_alpha[29][1] = 1'b1; \
	doodle_left_alpha[29][2] = 1'b1; \
	doodle_left_alpha[29][3] = 1'b1; \
	doodle_left_alpha[29][4] = 1'b1; \
	doodle_left_alpha[29][5] = 1'b1; \
	doodle_left_alpha[29][6] = 1'b1; \
	doodle_left_alpha[29][7] = 1'b1; \
	doodle_left_alpha[29][8] = 1'b1; \
	doodle_left_alpha[29][9] = 1'b1; \
	doodle_left_alpha[29][10] = 1'b1; \
	doodle_left_alpha[29][11] = 1'b1; \
	doodle_left_alpha[29][12] = 1'b1; \
	doodle_left_alpha[29][13] = 1'b1; \
	doodle_left_alpha[29][14] = 1'b1; \
	doodle_left_alpha[29][15] = 1'b1; \
	doodle_left_alpha[29][16] = 1'b1; \
	doodle_left_alpha[29][17] = 1'b1; \
	doodle_left_alpha[29][18] = 1'b1; \
	doodle_left_alpha[29][19] = 1'b1; \
	doodle_left_alpha[29][20] = 1'b1; \
	doodle_left_alpha[29][21] = 1'b1; \
	doodle_left_alpha[29][22] = 1'b1; \
	doodle_left_alpha[29][23] = 1'b0; \
	doodle_left_alpha[29][24] = 1'b0; \
	doodle_left_alpha[29][25] = 1'b0; \
	doodle_left_alpha[29][26] = 1'b0; \
	doodle_left_alpha[29][27] = 1'b0; \
	doodle_left_alpha[29][28] = 1'b0; \
	doodle_left_alpha[29][29] = 1'b0; \
	doodle_left_alpha[29][30] = 1'b0; \
	doodle_left_alpha[29][31] = 1'b0; \
	doodle_left_alpha[29][32] = 1'b0; \
	doodle_left_alpha[29][33] = 1'b0; \
	doodle_left_alpha[29][34] = 1'b0; \
	doodle_left_alpha[29][35] = 1'b0; \
	doodle_left_alpha[29][36] = 1'b0; \
	doodle_left_alpha[29][37] = 1'b0; \
	doodle_left_alpha[29][38] = 1'b0; \
	doodle_left_alpha[29][39] = 1'b0; \
	doodle_left_alpha[29][40] = 1'b0; \
	doodle_left_alpha[29][41] = 1'b0; \
	doodle_left_alpha[29][42] = 1'b0; \
	doodle_left_alpha[29][43] = 1'b0; \
	doodle_left_alpha[29][44] = 1'b0; \
	doodle_left_alpha[29][45] = 1'b0; \
	doodle_left_alpha[29][46] = 1'b0; \
	doodle_left_alpha[29][47] = 1'b0; \
	doodle_left_alpha[29][48] = 1'b0; \
	doodle_left_alpha[29][49] = 1'b0; \
	doodle_left_alpha[29][50] = 1'b0; \
	doodle_left_alpha[29][51] = 1'b0; \
	doodle_left_alpha[29][52] = 1'b0; \
	doodle_left_alpha[29][53] = 1'b0; \
	doodle_left_alpha[29][54] = 1'b0; \
	doodle_left_alpha[29][55] = 1'b0; \
	doodle_left_alpha[29][56] = 1'b0; \
	doodle_left_alpha[29][57] = 1'b0; \
	doodle_left_alpha[29][58] = 1'b0; \
	doodle_left_alpha[29][59] = 1'b0; \
	doodle_left_alpha[29][60] = 1'b0; \
	doodle_left_alpha[29][61] = 1'b0; \
	doodle_left_alpha[29][62] = 1'b0; \
	doodle_left_alpha[29][63] = 1'b0; \
	doodle_left_alpha[29][64] = 1'b0; \
	doodle_left_alpha[29][65] = 1'b1; \
	doodle_left_alpha[29][66] = 1'b1; \
	doodle_left_alpha[29][67] = 1'b1; \
	doodle_left_alpha[29][68] = 1'b1; \
	doodle_left_alpha[29][69] = 1'b1; \
	doodle_left_alpha[29][70] = 1'b1; \
	doodle_left_alpha[29][71] = 1'b1; \
	doodle_left_alpha[29][72] = 1'b1; \
	doodle_left_alpha[29][73] = 1'b1; \
	doodle_left_alpha[29][74] = 1'b1; \
	doodle_left_alpha[29][75] = 1'b1; \
	doodle_left_alpha[29][76] = 1'b1; \
	doodle_left_alpha[29][77] = 1'b1; \
	doodle_left_alpha[29][78] = 1'b1; \
	doodle_left_alpha[29][79] = 1'b1; \
	doodle_left_alpha[30][0] = 1'b1; \
	doodle_left_alpha[30][1] = 1'b1; \
	doodle_left_alpha[30][2] = 1'b1; \
	doodle_left_alpha[30][3] = 1'b1; \
	doodle_left_alpha[30][4] = 1'b1; \
	doodle_left_alpha[30][5] = 1'b1; \
	doodle_left_alpha[30][6] = 1'b1; \
	doodle_left_alpha[30][7] = 1'b1; \
	doodle_left_alpha[30][8] = 1'b1; \
	doodle_left_alpha[30][9] = 1'b1; \
	doodle_left_alpha[30][10] = 1'b1; \
	doodle_left_alpha[30][11] = 1'b1; \
	doodle_left_alpha[30][12] = 1'b1; \
	doodle_left_alpha[30][13] = 1'b1; \
	doodle_left_alpha[30][14] = 1'b1; \
	doodle_left_alpha[30][15] = 1'b1; \
	doodle_left_alpha[30][16] = 1'b1; \
	doodle_left_alpha[30][17] = 1'b1; \
	doodle_left_alpha[30][18] = 1'b1; \
	doodle_left_alpha[30][19] = 1'b1; \
	doodle_left_alpha[30][20] = 1'b1; \
	doodle_left_alpha[30][21] = 1'b1; \
	doodle_left_alpha[30][22] = 1'b1; \
	doodle_left_alpha[30][23] = 1'b0; \
	doodle_left_alpha[30][24] = 1'b0; \
	doodle_left_alpha[30][25] = 1'b0; \
	doodle_left_alpha[30][26] = 1'b0; \
	doodle_left_alpha[30][27] = 1'b0; \
	doodle_left_alpha[30][28] = 1'b0; \
	doodle_left_alpha[30][29] = 1'b0; \
	doodle_left_alpha[30][30] = 1'b0; \
	doodle_left_alpha[30][31] = 1'b0; \
	doodle_left_alpha[30][32] = 1'b0; \
	doodle_left_alpha[30][33] = 1'b0; \
	doodle_left_alpha[30][34] = 1'b0; \
	doodle_left_alpha[30][35] = 1'b0; \
	doodle_left_alpha[30][36] = 1'b0; \
	doodle_left_alpha[30][37] = 1'b0; \
	doodle_left_alpha[30][38] = 1'b0; \
	doodle_left_alpha[30][39] = 1'b0; \
	doodle_left_alpha[30][40] = 1'b0; \
	doodle_left_alpha[30][41] = 1'b0; \
	doodle_left_alpha[30][42] = 1'b0; \
	doodle_left_alpha[30][43] = 1'b0; \
	doodle_left_alpha[30][44] = 1'b0; \
	doodle_left_alpha[30][45] = 1'b0; \
	doodle_left_alpha[30][46] = 1'b0; \
	doodle_left_alpha[30][47] = 1'b0; \
	doodle_left_alpha[30][48] = 1'b0; \
	doodle_left_alpha[30][49] = 1'b0; \
	doodle_left_alpha[30][50] = 1'b0; \
	doodle_left_alpha[30][51] = 1'b0; \
	doodle_left_alpha[30][52] = 1'b0; \
	doodle_left_alpha[30][53] = 1'b0; \
	doodle_left_alpha[30][54] = 1'b0; \
	doodle_left_alpha[30][55] = 1'b0; \
	doodle_left_alpha[30][56] = 1'b0; \
	doodle_left_alpha[30][57] = 1'b0; \
	doodle_left_alpha[30][58] = 1'b0; \
	doodle_left_alpha[30][59] = 1'b0; \
	doodle_left_alpha[30][60] = 1'b0; \
	doodle_left_alpha[30][61] = 1'b0; \
	doodle_left_alpha[30][62] = 1'b0; \
	doodle_left_alpha[30][63] = 1'b0; \
	doodle_left_alpha[30][64] = 1'b0; \
	doodle_left_alpha[30][65] = 1'b1; \
	doodle_left_alpha[30][66] = 1'b1; \
	doodle_left_alpha[30][67] = 1'b1; \
	doodle_left_alpha[30][68] = 1'b1; \
	doodle_left_alpha[30][69] = 1'b1; \
	doodle_left_alpha[30][70] = 1'b1; \
	doodle_left_alpha[30][71] = 1'b1; \
	doodle_left_alpha[30][72] = 1'b1; \
	doodle_left_alpha[30][73] = 1'b1; \
	doodle_left_alpha[30][74] = 1'b1; \
	doodle_left_alpha[30][75] = 1'b1; \
	doodle_left_alpha[30][76] = 1'b1; \
	doodle_left_alpha[30][77] = 1'b1; \
	doodle_left_alpha[30][78] = 1'b1; \
	doodle_left_alpha[30][79] = 1'b1; \
	doodle_left_alpha[31][0] = 1'b1; \
	doodle_left_alpha[31][1] = 1'b1; \
	doodle_left_alpha[31][2] = 1'b1; \
	doodle_left_alpha[31][3] = 1'b1; \
	doodle_left_alpha[31][4] = 1'b1; \
	doodle_left_alpha[31][5] = 1'b1; \
	doodle_left_alpha[31][6] = 1'b1; \
	doodle_left_alpha[31][7] = 1'b1; \
	doodle_left_alpha[31][8] = 1'b1; \
	doodle_left_alpha[31][9] = 1'b1; \
	doodle_left_alpha[31][10] = 1'b1; \
	doodle_left_alpha[31][11] = 1'b1; \
	doodle_left_alpha[31][12] = 1'b1; \
	doodle_left_alpha[31][13] = 1'b1; \
	doodle_left_alpha[31][14] = 1'b1; \
	doodle_left_alpha[31][15] = 1'b1; \
	doodle_left_alpha[31][16] = 1'b1; \
	doodle_left_alpha[31][17] = 1'b1; \
	doodle_left_alpha[31][18] = 1'b1; \
	doodle_left_alpha[31][19] = 1'b1; \
	doodle_left_alpha[31][20] = 1'b1; \
	doodle_left_alpha[31][21] = 1'b1; \
	doodle_left_alpha[31][22] = 1'b1; \
	doodle_left_alpha[31][23] = 1'b0; \
	doodle_left_alpha[31][24] = 1'b0; \
	doodle_left_alpha[31][25] = 1'b0; \
	doodle_left_alpha[31][26] = 1'b0; \
	doodle_left_alpha[31][27] = 1'b0; \
	doodle_left_alpha[31][28] = 1'b0; \
	doodle_left_alpha[31][29] = 1'b0; \
	doodle_left_alpha[31][30] = 1'b0; \
	doodle_left_alpha[31][31] = 1'b0; \
	doodle_left_alpha[31][32] = 1'b0; \
	doodle_left_alpha[31][33] = 1'b0; \
	doodle_left_alpha[31][34] = 1'b0; \
	doodle_left_alpha[31][35] = 1'b0; \
	doodle_left_alpha[31][36] = 1'b0; \
	doodle_left_alpha[31][37] = 1'b0; \
	doodle_left_alpha[31][38] = 1'b0; \
	doodle_left_alpha[31][39] = 1'b0; \
	doodle_left_alpha[31][40] = 1'b0; \
	doodle_left_alpha[31][41] = 1'b0; \
	doodle_left_alpha[31][42] = 1'b0; \
	doodle_left_alpha[31][43] = 1'b0; \
	doodle_left_alpha[31][44] = 1'b0; \
	doodle_left_alpha[31][45] = 1'b0; \
	doodle_left_alpha[31][46] = 1'b0; \
	doodle_left_alpha[31][47] = 1'b0; \
	doodle_left_alpha[31][48] = 1'b0; \
	doodle_left_alpha[31][49] = 1'b0; \
	doodle_left_alpha[31][50] = 1'b0; \
	doodle_left_alpha[31][51] = 1'b0; \
	doodle_left_alpha[31][52] = 1'b0; \
	doodle_left_alpha[31][53] = 1'b0; \
	doodle_left_alpha[31][54] = 1'b0; \
	doodle_left_alpha[31][55] = 1'b0; \
	doodle_left_alpha[31][56] = 1'b0; \
	doodle_left_alpha[31][57] = 1'b0; \
	doodle_left_alpha[31][58] = 1'b0; \
	doodle_left_alpha[31][59] = 1'b0; \
	doodle_left_alpha[31][60] = 1'b0; \
	doodle_left_alpha[31][61] = 1'b0; \
	doodle_left_alpha[31][62] = 1'b0; \
	doodle_left_alpha[31][63] = 1'b0; \
	doodle_left_alpha[31][64] = 1'b0; \
	doodle_left_alpha[31][65] = 1'b1; \
	doodle_left_alpha[31][66] = 1'b1; \
	doodle_left_alpha[31][67] = 1'b1; \
	doodle_left_alpha[31][68] = 1'b1; \
	doodle_left_alpha[31][69] = 1'b1; \
	doodle_left_alpha[31][70] = 1'b1; \
	doodle_left_alpha[31][71] = 1'b1; \
	doodle_left_alpha[31][72] = 1'b1; \
	doodle_left_alpha[31][73] = 1'b1; \
	doodle_left_alpha[31][74] = 1'b1; \
	doodle_left_alpha[31][75] = 1'b1; \
	doodle_left_alpha[31][76] = 1'b1; \
	doodle_left_alpha[31][77] = 1'b1; \
	doodle_left_alpha[31][78] = 1'b1; \
	doodle_left_alpha[31][79] = 1'b1; \
	doodle_left_alpha[32][0] = 1'b1; \
	doodle_left_alpha[32][1] = 1'b1; \
	doodle_left_alpha[32][2] = 1'b1; \
	doodle_left_alpha[32][3] = 1'b1; \
	doodle_left_alpha[32][4] = 1'b1; \
	doodle_left_alpha[32][5] = 1'b1; \
	doodle_left_alpha[32][6] = 1'b1; \
	doodle_left_alpha[32][7] = 1'b1; \
	doodle_left_alpha[32][8] = 1'b1; \
	doodle_left_alpha[32][9] = 1'b1; \
	doodle_left_alpha[32][10] = 1'b1; \
	doodle_left_alpha[32][11] = 1'b1; \
	doodle_left_alpha[32][12] = 1'b1; \
	doodle_left_alpha[32][13] = 1'b1; \
	doodle_left_alpha[32][14] = 1'b1; \
	doodle_left_alpha[32][15] = 1'b1; \
	doodle_left_alpha[32][16] = 1'b1; \
	doodle_left_alpha[32][17] = 1'b1; \
	doodle_left_alpha[32][18] = 1'b1; \
	doodle_left_alpha[32][19] = 1'b1; \
	doodle_left_alpha[32][20] = 1'b1; \
	doodle_left_alpha[32][21] = 1'b1; \
	doodle_left_alpha[32][22] = 1'b1; \
	doodle_left_alpha[32][23] = 1'b0; \
	doodle_left_alpha[32][24] = 1'b0; \
	doodle_left_alpha[32][25] = 1'b0; \
	doodle_left_alpha[32][26] = 1'b0; \
	doodle_left_alpha[32][27] = 1'b0; \
	doodle_left_alpha[32][28] = 1'b0; \
	doodle_left_alpha[32][29] = 1'b0; \
	doodle_left_alpha[32][30] = 1'b0; \
	doodle_left_alpha[32][31] = 1'b0; \
	doodle_left_alpha[32][32] = 1'b0; \
	doodle_left_alpha[32][33] = 1'b0; \
	doodle_left_alpha[32][34] = 1'b0; \
	doodle_left_alpha[32][35] = 1'b0; \
	doodle_left_alpha[32][36] = 1'b0; \
	doodle_left_alpha[32][37] = 1'b0; \
	doodle_left_alpha[32][38] = 1'b0; \
	doodle_left_alpha[32][39] = 1'b0; \
	doodle_left_alpha[32][40] = 1'b0; \
	doodle_left_alpha[32][41] = 1'b0; \
	doodle_left_alpha[32][42] = 1'b0; \
	doodle_left_alpha[32][43] = 1'b0; \
	doodle_left_alpha[32][44] = 1'b0; \
	doodle_left_alpha[32][45] = 1'b0; \
	doodle_left_alpha[32][46] = 1'b0; \
	doodle_left_alpha[32][47] = 1'b0; \
	doodle_left_alpha[32][48] = 1'b0; \
	doodle_left_alpha[32][49] = 1'b0; \
	doodle_left_alpha[32][50] = 1'b0; \
	doodle_left_alpha[32][51] = 1'b0; \
	doodle_left_alpha[32][52] = 1'b0; \
	doodle_left_alpha[32][53] = 1'b0; \
	doodle_left_alpha[32][54] = 1'b0; \
	doodle_left_alpha[32][55] = 1'b0; \
	doodle_left_alpha[32][56] = 1'b0; \
	doodle_left_alpha[32][57] = 1'b0; \
	doodle_left_alpha[32][58] = 1'b0; \
	doodle_left_alpha[32][59] = 1'b0; \
	doodle_left_alpha[32][60] = 1'b0; \
	doodle_left_alpha[32][61] = 1'b0; \
	doodle_left_alpha[32][62] = 1'b0; \
	doodle_left_alpha[32][63] = 1'b0; \
	doodle_left_alpha[32][64] = 1'b0; \
	doodle_left_alpha[32][65] = 1'b1; \
	doodle_left_alpha[32][66] = 1'b1; \
	doodle_left_alpha[32][67] = 1'b1; \
	doodle_left_alpha[32][68] = 1'b1; \
	doodle_left_alpha[32][69] = 1'b1; \
	doodle_left_alpha[32][70] = 1'b1; \
	doodle_left_alpha[32][71] = 1'b1; \
	doodle_left_alpha[32][72] = 1'b1; \
	doodle_left_alpha[32][73] = 1'b1; \
	doodle_left_alpha[32][74] = 1'b1; \
	doodle_left_alpha[32][75] = 1'b1; \
	doodle_left_alpha[32][76] = 1'b1; \
	doodle_left_alpha[32][77] = 1'b1; \
	doodle_left_alpha[32][78] = 1'b1; \
	doodle_left_alpha[32][79] = 1'b1; \
	doodle_left_alpha[33][0] = 1'b1; \
	doodle_left_alpha[33][1] = 1'b1; \
	doodle_left_alpha[33][2] = 1'b1; \
	doodle_left_alpha[33][3] = 1'b1; \
	doodle_left_alpha[33][4] = 1'b1; \
	doodle_left_alpha[33][5] = 1'b1; \
	doodle_left_alpha[33][6] = 1'b1; \
	doodle_left_alpha[33][7] = 1'b1; \
	doodle_left_alpha[33][8] = 1'b1; \
	doodle_left_alpha[33][9] = 1'b1; \
	doodle_left_alpha[33][10] = 1'b1; \
	doodle_left_alpha[33][11] = 1'b1; \
	doodle_left_alpha[33][12] = 1'b1; \
	doodle_left_alpha[33][13] = 1'b1; \
	doodle_left_alpha[33][14] = 1'b1; \
	doodle_left_alpha[33][15] = 1'b1; \
	doodle_left_alpha[33][16] = 1'b1; \
	doodle_left_alpha[33][17] = 1'b1; \
	doodle_left_alpha[33][18] = 1'b1; \
	doodle_left_alpha[33][19] = 1'b1; \
	doodle_left_alpha[33][20] = 1'b1; \
	doodle_left_alpha[33][21] = 1'b1; \
	doodle_left_alpha[33][22] = 1'b1; \
	doodle_left_alpha[33][23] = 1'b0; \
	doodle_left_alpha[33][24] = 1'b0; \
	doodle_left_alpha[33][25] = 1'b0; \
	doodle_left_alpha[33][26] = 1'b0; \
	doodle_left_alpha[33][27] = 1'b0; \
	doodle_left_alpha[33][28] = 1'b0; \
	doodle_left_alpha[33][29] = 1'b0; \
	doodle_left_alpha[33][30] = 1'b0; \
	doodle_left_alpha[33][31] = 1'b0; \
	doodle_left_alpha[33][32] = 1'b0; \
	doodle_left_alpha[33][33] = 1'b0; \
	doodle_left_alpha[33][34] = 1'b0; \
	doodle_left_alpha[33][35] = 1'b0; \
	doodle_left_alpha[33][36] = 1'b0; \
	doodle_left_alpha[33][37] = 1'b0; \
	doodle_left_alpha[33][38] = 1'b0; \
	doodle_left_alpha[33][39] = 1'b0; \
	doodle_left_alpha[33][40] = 1'b0; \
	doodle_left_alpha[33][41] = 1'b0; \
	doodle_left_alpha[33][42] = 1'b0; \
	doodle_left_alpha[33][43] = 1'b0; \
	doodle_left_alpha[33][44] = 1'b0; \
	doodle_left_alpha[33][45] = 1'b0; \
	doodle_left_alpha[33][46] = 1'b0; \
	doodle_left_alpha[33][47] = 1'b0; \
	doodle_left_alpha[33][48] = 1'b0; \
	doodle_left_alpha[33][49] = 1'b0; \
	doodle_left_alpha[33][50] = 1'b0; \
	doodle_left_alpha[33][51] = 1'b0; \
	doodle_left_alpha[33][52] = 1'b0; \
	doodle_left_alpha[33][53] = 1'b0; \
	doodle_left_alpha[33][54] = 1'b0; \
	doodle_left_alpha[33][55] = 1'b0; \
	doodle_left_alpha[33][56] = 1'b0; \
	doodle_left_alpha[33][57] = 1'b0; \
	doodle_left_alpha[33][58] = 1'b0; \
	doodle_left_alpha[33][59] = 1'b0; \
	doodle_left_alpha[33][60] = 1'b0; \
	doodle_left_alpha[33][61] = 1'b0; \
	doodle_left_alpha[33][62] = 1'b0; \
	doodle_left_alpha[33][63] = 1'b0; \
	doodle_left_alpha[33][64] = 1'b0; \
	doodle_left_alpha[33][65] = 1'b1; \
	doodle_left_alpha[33][66] = 1'b1; \
	doodle_left_alpha[33][67] = 1'b1; \
	doodle_left_alpha[33][68] = 1'b1; \
	doodle_left_alpha[33][69] = 1'b1; \
	doodle_left_alpha[33][70] = 1'b1; \
	doodle_left_alpha[33][71] = 1'b1; \
	doodle_left_alpha[33][72] = 1'b1; \
	doodle_left_alpha[33][73] = 1'b1; \
	doodle_left_alpha[33][74] = 1'b1; \
	doodle_left_alpha[33][75] = 1'b1; \
	doodle_left_alpha[33][76] = 1'b1; \
	doodle_left_alpha[33][77] = 1'b1; \
	doodle_left_alpha[33][78] = 1'b1; \
	doodle_left_alpha[33][79] = 1'b1; \
	doodle_left_alpha[34][0] = 1'b1; \
	doodle_left_alpha[34][1] = 1'b1; \
	doodle_left_alpha[34][2] = 1'b1; \
	doodle_left_alpha[34][3] = 1'b1; \
	doodle_left_alpha[34][4] = 1'b0; \
	doodle_left_alpha[34][5] = 1'b0; \
	doodle_left_alpha[34][6] = 1'b0; \
	doodle_left_alpha[34][7] = 1'b0; \
	doodle_left_alpha[34][8] = 1'b0; \
	doodle_left_alpha[34][9] = 1'b0; \
	doodle_left_alpha[34][10] = 1'b0; \
	doodle_left_alpha[34][11] = 1'b0; \
	doodle_left_alpha[34][12] = 1'b0; \
	doodle_left_alpha[34][13] = 1'b0; \
	doodle_left_alpha[34][14] = 1'b0; \
	doodle_left_alpha[34][15] = 1'b0; \
	doodle_left_alpha[34][16] = 1'b0; \
	doodle_left_alpha[34][17] = 1'b0; \
	doodle_left_alpha[34][18] = 1'b0; \
	doodle_left_alpha[34][19] = 1'b0; \
	doodle_left_alpha[34][20] = 1'b0; \
	doodle_left_alpha[34][21] = 1'b0; \
	doodle_left_alpha[34][22] = 1'b0; \
	doodle_left_alpha[34][23] = 1'b0; \
	doodle_left_alpha[34][24] = 1'b0; \
	doodle_left_alpha[34][25] = 1'b0; \
	doodle_left_alpha[34][26] = 1'b0; \
	doodle_left_alpha[34][27] = 1'b0; \
	doodle_left_alpha[34][28] = 1'b0; \
	doodle_left_alpha[34][29] = 1'b0; \
	doodle_left_alpha[34][30] = 1'b0; \
	doodle_left_alpha[34][31] = 1'b0; \
	doodle_left_alpha[34][32] = 1'b0; \
	doodle_left_alpha[34][33] = 1'b0; \
	doodle_left_alpha[34][34] = 1'b0; \
	doodle_left_alpha[34][35] = 1'b0; \
	doodle_left_alpha[34][36] = 1'b0; \
	doodle_left_alpha[34][37] = 1'b0; \
	doodle_left_alpha[34][38] = 1'b0; \
	doodle_left_alpha[34][39] = 1'b0; \
	doodle_left_alpha[34][40] = 1'b0; \
	doodle_left_alpha[34][41] = 1'b0; \
	doodle_left_alpha[34][42] = 1'b0; \
	doodle_left_alpha[34][43] = 1'b0; \
	doodle_left_alpha[34][44] = 1'b0; \
	doodle_left_alpha[34][45] = 1'b0; \
	doodle_left_alpha[34][46] = 1'b0; \
	doodle_left_alpha[34][47] = 1'b0; \
	doodle_left_alpha[34][48] = 1'b0; \
	doodle_left_alpha[34][49] = 1'b0; \
	doodle_left_alpha[34][50] = 1'b0; \
	doodle_left_alpha[34][51] = 1'b0; \
	doodle_left_alpha[34][52] = 1'b0; \
	doodle_left_alpha[34][53] = 1'b0; \
	doodle_left_alpha[34][54] = 1'b0; \
	doodle_left_alpha[34][55] = 1'b0; \
	doodle_left_alpha[34][56] = 1'b0; \
	doodle_left_alpha[34][57] = 1'b0; \
	doodle_left_alpha[34][58] = 1'b0; \
	doodle_left_alpha[34][59] = 1'b0; \
	doodle_left_alpha[34][60] = 1'b0; \
	doodle_left_alpha[34][61] = 1'b0; \
	doodle_left_alpha[34][62] = 1'b0; \
	doodle_left_alpha[34][63] = 1'b0; \
	doodle_left_alpha[34][64] = 1'b0; \
	doodle_left_alpha[34][65] = 1'b1; \
	doodle_left_alpha[34][66] = 1'b1; \
	doodle_left_alpha[34][67] = 1'b1; \
	doodle_left_alpha[34][68] = 1'b1; \
	doodle_left_alpha[34][69] = 1'b1; \
	doodle_left_alpha[34][70] = 1'b1; \
	doodle_left_alpha[34][71] = 1'b1; \
	doodle_left_alpha[34][72] = 1'b1; \
	doodle_left_alpha[34][73] = 1'b1; \
	doodle_left_alpha[34][74] = 1'b1; \
	doodle_left_alpha[34][75] = 1'b1; \
	doodle_left_alpha[34][76] = 1'b1; \
	doodle_left_alpha[34][77] = 1'b1; \
	doodle_left_alpha[34][78] = 1'b1; \
	doodle_left_alpha[34][79] = 1'b1; \
	doodle_left_alpha[35][0] = 1'b1; \
	doodle_left_alpha[35][1] = 1'b1; \
	doodle_left_alpha[35][2] = 1'b1; \
	doodle_left_alpha[35][3] = 1'b1; \
	doodle_left_alpha[35][4] = 1'b0; \
	doodle_left_alpha[35][5] = 1'b0; \
	doodle_left_alpha[35][6] = 1'b0; \
	doodle_left_alpha[35][7] = 1'b0; \
	doodle_left_alpha[35][8] = 1'b0; \
	doodle_left_alpha[35][9] = 1'b0; \
	doodle_left_alpha[35][10] = 1'b0; \
	doodle_left_alpha[35][11] = 1'b0; \
	doodle_left_alpha[35][12] = 1'b0; \
	doodle_left_alpha[35][13] = 1'b0; \
	doodle_left_alpha[35][14] = 1'b0; \
	doodle_left_alpha[35][15] = 1'b0; \
	doodle_left_alpha[35][16] = 1'b0; \
	doodle_left_alpha[35][17] = 1'b0; \
	doodle_left_alpha[35][18] = 1'b0; \
	doodle_left_alpha[35][19] = 1'b0; \
	doodle_left_alpha[35][20] = 1'b0; \
	doodle_left_alpha[35][21] = 1'b0; \
	doodle_left_alpha[35][22] = 1'b0; \
	doodle_left_alpha[35][23] = 1'b0; \
	doodle_left_alpha[35][24] = 1'b0; \
	doodle_left_alpha[35][25] = 1'b0; \
	doodle_left_alpha[35][26] = 1'b0; \
	doodle_left_alpha[35][27] = 1'b0; \
	doodle_left_alpha[35][28] = 1'b0; \
	doodle_left_alpha[35][29] = 1'b0; \
	doodle_left_alpha[35][30] = 1'b0; \
	doodle_left_alpha[35][31] = 1'b0; \
	doodle_left_alpha[35][32] = 1'b0; \
	doodle_left_alpha[35][33] = 1'b0; \
	doodle_left_alpha[35][34] = 1'b0; \
	doodle_left_alpha[35][35] = 1'b0; \
	doodle_left_alpha[35][36] = 1'b0; \
	doodle_left_alpha[35][37] = 1'b0; \
	doodle_left_alpha[35][38] = 1'b0; \
	doodle_left_alpha[35][39] = 1'b0; \
	doodle_left_alpha[35][40] = 1'b0; \
	doodle_left_alpha[35][41] = 1'b0; \
	doodle_left_alpha[35][42] = 1'b0; \
	doodle_left_alpha[35][43] = 1'b0; \
	doodle_left_alpha[35][44] = 1'b0; \
	doodle_left_alpha[35][45] = 1'b0; \
	doodle_left_alpha[35][46] = 1'b0; \
	doodle_left_alpha[35][47] = 1'b0; \
	doodle_left_alpha[35][48] = 1'b0; \
	doodle_left_alpha[35][49] = 1'b0; \
	doodle_left_alpha[35][50] = 1'b0; \
	doodle_left_alpha[35][51] = 1'b0; \
	doodle_left_alpha[35][52] = 1'b0; \
	doodle_left_alpha[35][53] = 1'b0; \
	doodle_left_alpha[35][54] = 1'b0; \
	doodle_left_alpha[35][55] = 1'b0; \
	doodle_left_alpha[35][56] = 1'b0; \
	doodle_left_alpha[35][57] = 1'b0; \
	doodle_left_alpha[35][58] = 1'b0; \
	doodle_left_alpha[35][59] = 1'b0; \
	doodle_left_alpha[35][60] = 1'b0; \
	doodle_left_alpha[35][61] = 1'b0; \
	doodle_left_alpha[35][62] = 1'b0; \
	doodle_left_alpha[35][63] = 1'b0; \
	doodle_left_alpha[35][64] = 1'b0; \
	doodle_left_alpha[35][65] = 1'b1; \
	doodle_left_alpha[35][66] = 1'b1; \
	doodle_left_alpha[35][67] = 1'b1; \
	doodle_left_alpha[35][68] = 1'b1; \
	doodle_left_alpha[35][69] = 1'b1; \
	doodle_left_alpha[35][70] = 1'b1; \
	doodle_left_alpha[35][71] = 1'b1; \
	doodle_left_alpha[35][72] = 1'b1; \
	doodle_left_alpha[35][73] = 1'b1; \
	doodle_left_alpha[35][74] = 1'b1; \
	doodle_left_alpha[35][75] = 1'b1; \
	doodle_left_alpha[35][76] = 1'b1; \
	doodle_left_alpha[35][77] = 1'b1; \
	doodle_left_alpha[35][78] = 1'b1; \
	doodle_left_alpha[35][79] = 1'b1; \
	doodle_left_alpha[36][0] = 1'b1; \
	doodle_left_alpha[36][1] = 1'b1; \
	doodle_left_alpha[36][2] = 1'b1; \
	doodle_left_alpha[36][3] = 1'b1; \
	doodle_left_alpha[36][4] = 1'b0; \
	doodle_left_alpha[36][5] = 1'b0; \
	doodle_left_alpha[36][6] = 1'b0; \
	doodle_left_alpha[36][7] = 1'b0; \
	doodle_left_alpha[36][8] = 1'b0; \
	doodle_left_alpha[36][9] = 1'b0; \
	doodle_left_alpha[36][10] = 1'b0; \
	doodle_left_alpha[36][11] = 1'b0; \
	doodle_left_alpha[36][12] = 1'b0; \
	doodle_left_alpha[36][13] = 1'b0; \
	doodle_left_alpha[36][14] = 1'b0; \
	doodle_left_alpha[36][15] = 1'b0; \
	doodle_left_alpha[36][16] = 1'b0; \
	doodle_left_alpha[36][17] = 1'b0; \
	doodle_left_alpha[36][18] = 1'b0; \
	doodle_left_alpha[36][19] = 1'b0; \
	doodle_left_alpha[36][20] = 1'b0; \
	doodle_left_alpha[36][21] = 1'b0; \
	doodle_left_alpha[36][22] = 1'b0; \
	doodle_left_alpha[36][23] = 1'b0; \
	doodle_left_alpha[36][24] = 1'b0; \
	doodle_left_alpha[36][25] = 1'b0; \
	doodle_left_alpha[36][26] = 1'b0; \
	doodle_left_alpha[36][27] = 1'b0; \
	doodle_left_alpha[36][28] = 1'b0; \
	doodle_left_alpha[36][29] = 1'b0; \
	doodle_left_alpha[36][30] = 1'b0; \
	doodle_left_alpha[36][31] = 1'b0; \
	doodle_left_alpha[36][32] = 1'b0; \
	doodle_left_alpha[36][33] = 1'b0; \
	doodle_left_alpha[36][34] = 1'b0; \
	doodle_left_alpha[36][35] = 1'b0; \
	doodle_left_alpha[36][36] = 1'b0; \
	doodle_left_alpha[36][37] = 1'b0; \
	doodle_left_alpha[36][38] = 1'b0; \
	doodle_left_alpha[36][39] = 1'b0; \
	doodle_left_alpha[36][40] = 1'b0; \
	doodle_left_alpha[36][41] = 1'b0; \
	doodle_left_alpha[36][42] = 1'b0; \
	doodle_left_alpha[36][43] = 1'b0; \
	doodle_left_alpha[36][44] = 1'b0; \
	doodle_left_alpha[36][45] = 1'b0; \
	doodle_left_alpha[36][46] = 1'b0; \
	doodle_left_alpha[36][47] = 1'b0; \
	doodle_left_alpha[36][48] = 1'b0; \
	doodle_left_alpha[36][49] = 1'b0; \
	doodle_left_alpha[36][50] = 1'b0; \
	doodle_left_alpha[36][51] = 1'b0; \
	doodle_left_alpha[36][52] = 1'b0; \
	doodle_left_alpha[36][53] = 1'b0; \
	doodle_left_alpha[36][54] = 1'b0; \
	doodle_left_alpha[36][55] = 1'b0; \
	doodle_left_alpha[36][56] = 1'b0; \
	doodle_left_alpha[36][57] = 1'b0; \
	doodle_left_alpha[36][58] = 1'b0; \
	doodle_left_alpha[36][59] = 1'b0; \
	doodle_left_alpha[36][60] = 1'b0; \
	doodle_left_alpha[36][61] = 1'b0; \
	doodle_left_alpha[36][62] = 1'b0; \
	doodle_left_alpha[36][63] = 1'b0; \
	doodle_left_alpha[36][64] = 1'b0; \
	doodle_left_alpha[36][65] = 1'b1; \
	doodle_left_alpha[36][66] = 1'b1; \
	doodle_left_alpha[36][67] = 1'b1; \
	doodle_left_alpha[36][68] = 1'b1; \
	doodle_left_alpha[36][69] = 1'b1; \
	doodle_left_alpha[36][70] = 1'b1; \
	doodle_left_alpha[36][71] = 1'b1; \
	doodle_left_alpha[36][72] = 1'b1; \
	doodle_left_alpha[36][73] = 1'b1; \
	doodle_left_alpha[36][74] = 1'b1; \
	doodle_left_alpha[36][75] = 1'b1; \
	doodle_left_alpha[36][76] = 1'b1; \
	doodle_left_alpha[36][77] = 1'b1; \
	doodle_left_alpha[36][78] = 1'b1; \
	doodle_left_alpha[36][79] = 1'b1; \
	doodle_left_alpha[37][0] = 1'b1; \
	doodle_left_alpha[37][1] = 1'b1; \
	doodle_left_alpha[37][2] = 1'b1; \
	doodle_left_alpha[37][3] = 1'b1; \
	doodle_left_alpha[37][4] = 1'b0; \
	doodle_left_alpha[37][5] = 1'b0; \
	doodle_left_alpha[37][6] = 1'b0; \
	doodle_left_alpha[37][7] = 1'b0; \
	doodle_left_alpha[37][8] = 1'b0; \
	doodle_left_alpha[37][9] = 1'b0; \
	doodle_left_alpha[37][10] = 1'b0; \
	doodle_left_alpha[37][11] = 1'b0; \
	doodle_left_alpha[37][12] = 1'b0; \
	doodle_left_alpha[37][13] = 1'b0; \
	doodle_left_alpha[37][14] = 1'b0; \
	doodle_left_alpha[37][15] = 1'b0; \
	doodle_left_alpha[37][16] = 1'b0; \
	doodle_left_alpha[37][17] = 1'b0; \
	doodle_left_alpha[37][18] = 1'b0; \
	doodle_left_alpha[37][19] = 1'b0; \
	doodle_left_alpha[37][20] = 1'b0; \
	doodle_left_alpha[37][21] = 1'b0; \
	doodle_left_alpha[37][22] = 1'b0; \
	doodle_left_alpha[37][23] = 1'b0; \
	doodle_left_alpha[37][24] = 1'b0; \
	doodle_left_alpha[37][25] = 1'b0; \
	doodle_left_alpha[37][26] = 1'b0; \
	doodle_left_alpha[37][27] = 1'b0; \
	doodle_left_alpha[37][28] = 1'b0; \
	doodle_left_alpha[37][29] = 1'b0; \
	doodle_left_alpha[37][30] = 1'b0; \
	doodle_left_alpha[37][31] = 1'b0; \
	doodle_left_alpha[37][32] = 1'b0; \
	doodle_left_alpha[37][33] = 1'b0; \
	doodle_left_alpha[37][34] = 1'b0; \
	doodle_left_alpha[37][35] = 1'b0; \
	doodle_left_alpha[37][36] = 1'b0; \
	doodle_left_alpha[37][37] = 1'b0; \
	doodle_left_alpha[37][38] = 1'b0; \
	doodle_left_alpha[37][39] = 1'b0; \
	doodle_left_alpha[37][40] = 1'b0; \
	doodle_left_alpha[37][41] = 1'b0; \
	doodle_left_alpha[37][42] = 1'b0; \
	doodle_left_alpha[37][43] = 1'b0; \
	doodle_left_alpha[37][44] = 1'b0; \
	doodle_left_alpha[37][45] = 1'b0; \
	doodle_left_alpha[37][46] = 1'b0; \
	doodle_left_alpha[37][47] = 1'b0; \
	doodle_left_alpha[37][48] = 1'b0; \
	doodle_left_alpha[37][49] = 1'b0; \
	doodle_left_alpha[37][50] = 1'b0; \
	doodle_left_alpha[37][51] = 1'b0; \
	doodle_left_alpha[37][52] = 1'b0; \
	doodle_left_alpha[37][53] = 1'b0; \
	doodle_left_alpha[37][54] = 1'b0; \
	doodle_left_alpha[37][55] = 1'b0; \
	doodle_left_alpha[37][56] = 1'b0; \
	doodle_left_alpha[37][57] = 1'b0; \
	doodle_left_alpha[37][58] = 1'b0; \
	doodle_left_alpha[37][59] = 1'b0; \
	doodle_left_alpha[37][60] = 1'b0; \
	doodle_left_alpha[37][61] = 1'b0; \
	doodle_left_alpha[37][62] = 1'b0; \
	doodle_left_alpha[37][63] = 1'b0; \
	doodle_left_alpha[37][64] = 1'b0; \
	doodle_left_alpha[37][65] = 1'b1; \
	doodle_left_alpha[37][66] = 1'b1; \
	doodle_left_alpha[37][67] = 1'b1; \
	doodle_left_alpha[37][68] = 1'b1; \
	doodle_left_alpha[37][69] = 1'b1; \
	doodle_left_alpha[37][70] = 1'b1; \
	doodle_left_alpha[37][71] = 1'b1; \
	doodle_left_alpha[37][72] = 1'b1; \
	doodle_left_alpha[37][73] = 1'b1; \
	doodle_left_alpha[37][74] = 1'b1; \
	doodle_left_alpha[37][75] = 1'b1; \
	doodle_left_alpha[37][76] = 1'b1; \
	doodle_left_alpha[37][77] = 1'b1; \
	doodle_left_alpha[37][78] = 1'b1; \
	doodle_left_alpha[37][79] = 1'b1; \
	doodle_left_alpha[38][0] = 1'b1; \
	doodle_left_alpha[38][1] = 1'b1; \
	doodle_left_alpha[38][2] = 1'b1; \
	doodle_left_alpha[38][3] = 1'b1; \
	doodle_left_alpha[38][4] = 1'b0; \
	doodle_left_alpha[38][5] = 1'b0; \
	doodle_left_alpha[38][6] = 1'b0; \
	doodle_left_alpha[38][7] = 1'b0; \
	doodle_left_alpha[38][8] = 1'b0; \
	doodle_left_alpha[38][9] = 1'b0; \
	doodle_left_alpha[38][10] = 1'b0; \
	doodle_left_alpha[38][11] = 1'b0; \
	doodle_left_alpha[38][12] = 1'b0; \
	doodle_left_alpha[38][13] = 1'b0; \
	doodle_left_alpha[38][14] = 1'b0; \
	doodle_left_alpha[38][15] = 1'b0; \
	doodle_left_alpha[38][16] = 1'b0; \
	doodle_left_alpha[38][17] = 1'b0; \
	doodle_left_alpha[38][18] = 1'b0; \
	doodle_left_alpha[38][19] = 1'b0; \
	doodle_left_alpha[38][20] = 1'b0; \
	doodle_left_alpha[38][21] = 1'b0; \
	doodle_left_alpha[38][22] = 1'b0; \
	doodle_left_alpha[38][23] = 1'b0; \
	doodle_left_alpha[38][24] = 1'b0; \
	doodle_left_alpha[38][25] = 1'b0; \
	doodle_left_alpha[38][26] = 1'b0; \
	doodle_left_alpha[38][27] = 1'b0; \
	doodle_left_alpha[38][28] = 1'b0; \
	doodle_left_alpha[38][29] = 1'b0; \
	doodle_left_alpha[38][30] = 1'b0; \
	doodle_left_alpha[38][31] = 1'b0; \
	doodle_left_alpha[38][32] = 1'b0; \
	doodle_left_alpha[38][33] = 1'b0; \
	doodle_left_alpha[38][34] = 1'b0; \
	doodle_left_alpha[38][35] = 1'b0; \
	doodle_left_alpha[38][36] = 1'b0; \
	doodle_left_alpha[38][37] = 1'b0; \
	doodle_left_alpha[38][38] = 1'b0; \
	doodle_left_alpha[38][39] = 1'b0; \
	doodle_left_alpha[38][40] = 1'b0; \
	doodle_left_alpha[38][41] = 1'b0; \
	doodle_left_alpha[38][42] = 1'b0; \
	doodle_left_alpha[38][43] = 1'b0; \
	doodle_left_alpha[38][44] = 1'b0; \
	doodle_left_alpha[38][45] = 1'b0; \
	doodle_left_alpha[38][46] = 1'b0; \
	doodle_left_alpha[38][47] = 1'b0; \
	doodle_left_alpha[38][48] = 1'b0; \
	doodle_left_alpha[38][49] = 1'b0; \
	doodle_left_alpha[38][50] = 1'b0; \
	doodle_left_alpha[38][51] = 1'b0; \
	doodle_left_alpha[38][52] = 1'b0; \
	doodle_left_alpha[38][53] = 1'b0; \
	doodle_left_alpha[38][54] = 1'b0; \
	doodle_left_alpha[38][55] = 1'b0; \
	doodle_left_alpha[38][56] = 1'b0; \
	doodle_left_alpha[38][57] = 1'b0; \
	doodle_left_alpha[38][58] = 1'b0; \
	doodle_left_alpha[38][59] = 1'b0; \
	doodle_left_alpha[38][60] = 1'b0; \
	doodle_left_alpha[38][61] = 1'b0; \
	doodle_left_alpha[38][62] = 1'b0; \
	doodle_left_alpha[38][63] = 1'b0; \
	doodle_left_alpha[38][64] = 1'b0; \
	doodle_left_alpha[38][65] = 1'b1; \
	doodle_left_alpha[38][66] = 1'b1; \
	doodle_left_alpha[38][67] = 1'b1; \
	doodle_left_alpha[38][68] = 1'b1; \
	doodle_left_alpha[38][69] = 1'b1; \
	doodle_left_alpha[38][70] = 1'b1; \
	doodle_left_alpha[38][71] = 1'b1; \
	doodle_left_alpha[38][72] = 1'b1; \
	doodle_left_alpha[38][73] = 1'b1; \
	doodle_left_alpha[38][74] = 1'b1; \
	doodle_left_alpha[38][75] = 1'b1; \
	doodle_left_alpha[38][76] = 1'b1; \
	doodle_left_alpha[38][77] = 1'b1; \
	doodle_left_alpha[38][78] = 1'b1; \
	doodle_left_alpha[38][79] = 1'b1; \
	doodle_left_alpha[39][0] = 1'b1; \
	doodle_left_alpha[39][1] = 1'b1; \
	doodle_left_alpha[39][2] = 1'b1; \
	doodle_left_alpha[39][3] = 1'b1; \
	doodle_left_alpha[39][4] = 1'b0; \
	doodle_left_alpha[39][5] = 1'b0; \
	doodle_left_alpha[39][6] = 1'b0; \
	doodle_left_alpha[39][7] = 1'b0; \
	doodle_left_alpha[39][8] = 1'b0; \
	doodle_left_alpha[39][9] = 1'b0; \
	doodle_left_alpha[39][10] = 1'b0; \
	doodle_left_alpha[39][11] = 1'b0; \
	doodle_left_alpha[39][12] = 1'b0; \
	doodle_left_alpha[39][13] = 1'b0; \
	doodle_left_alpha[39][14] = 1'b0; \
	doodle_left_alpha[39][15] = 1'b0; \
	doodle_left_alpha[39][16] = 1'b0; \
	doodle_left_alpha[39][17] = 1'b0; \
	doodle_left_alpha[39][18] = 1'b0; \
	doodle_left_alpha[39][19] = 1'b0; \
	doodle_left_alpha[39][20] = 1'b0; \
	doodle_left_alpha[39][21] = 1'b0; \
	doodle_left_alpha[39][22] = 1'b0; \
	doodle_left_alpha[39][23] = 1'b0; \
	doodle_left_alpha[39][24] = 1'b0; \
	doodle_left_alpha[39][25] = 1'b0; \
	doodle_left_alpha[39][26] = 1'b0; \
	doodle_left_alpha[39][27] = 1'b0; \
	doodle_left_alpha[39][28] = 1'b0; \
	doodle_left_alpha[39][29] = 1'b0; \
	doodle_left_alpha[39][30] = 1'b0; \
	doodle_left_alpha[39][31] = 1'b0; \
	doodle_left_alpha[39][32] = 1'b0; \
	doodle_left_alpha[39][33] = 1'b0; \
	doodle_left_alpha[39][34] = 1'b0; \
	doodle_left_alpha[39][35] = 1'b0; \
	doodle_left_alpha[39][36] = 1'b0; \
	doodle_left_alpha[39][37] = 1'b0; \
	doodle_left_alpha[39][38] = 1'b0; \
	doodle_left_alpha[39][39] = 1'b0; \
	doodle_left_alpha[39][40] = 1'b0; \
	doodle_left_alpha[39][41] = 1'b0; \
	doodle_left_alpha[39][42] = 1'b0; \
	doodle_left_alpha[39][43] = 1'b0; \
	doodle_left_alpha[39][44] = 1'b0; \
	doodle_left_alpha[39][45] = 1'b0; \
	doodle_left_alpha[39][46] = 1'b0; \
	doodle_left_alpha[39][47] = 1'b0; \
	doodle_left_alpha[39][48] = 1'b0; \
	doodle_left_alpha[39][49] = 1'b0; \
	doodle_left_alpha[39][50] = 1'b0; \
	doodle_left_alpha[39][51] = 1'b0; \
	doodle_left_alpha[39][52] = 1'b0; \
	doodle_left_alpha[39][53] = 1'b0; \
	doodle_left_alpha[39][54] = 1'b0; \
	doodle_left_alpha[39][55] = 1'b0; \
	doodle_left_alpha[39][56] = 1'b0; \
	doodle_left_alpha[39][57] = 1'b0; \
	doodle_left_alpha[39][58] = 1'b0; \
	doodle_left_alpha[39][59] = 1'b0; \
	doodle_left_alpha[39][60] = 1'b0; \
	doodle_left_alpha[39][61] = 1'b0; \
	doodle_left_alpha[39][62] = 1'b0; \
	doodle_left_alpha[39][63] = 1'b0; \
	doodle_left_alpha[39][64] = 1'b0; \
	doodle_left_alpha[39][65] = 1'b1; \
	doodle_left_alpha[39][66] = 1'b1; \
	doodle_left_alpha[39][67] = 1'b1; \
	doodle_left_alpha[39][68] = 1'b1; \
	doodle_left_alpha[39][69] = 1'b1; \
	doodle_left_alpha[39][70] = 1'b1; \
	doodle_left_alpha[39][71] = 1'b1; \
	doodle_left_alpha[39][72] = 1'b1; \
	doodle_left_alpha[39][73] = 1'b1; \
	doodle_left_alpha[39][74] = 1'b1; \
	doodle_left_alpha[39][75] = 1'b1; \
	doodle_left_alpha[39][76] = 1'b1; \
	doodle_left_alpha[39][77] = 1'b1; \
	doodle_left_alpha[39][78] = 1'b1; \
	doodle_left_alpha[39][79] = 1'b1; \
	doodle_left_alpha[40][0] = 1'b1; \
	doodle_left_alpha[40][1] = 1'b1; \
	doodle_left_alpha[40][2] = 1'b1; \
	doodle_left_alpha[40][3] = 1'b1; \
	doodle_left_alpha[40][4] = 1'b0; \
	doodle_left_alpha[40][5] = 1'b0; \
	doodle_left_alpha[40][6] = 1'b0; \
	doodle_left_alpha[40][7] = 1'b0; \
	doodle_left_alpha[40][8] = 1'b0; \
	doodle_left_alpha[40][9] = 1'b0; \
	doodle_left_alpha[40][10] = 1'b0; \
	doodle_left_alpha[40][11] = 1'b0; \
	doodle_left_alpha[40][12] = 1'b0; \
	doodle_left_alpha[40][13] = 1'b0; \
	doodle_left_alpha[40][14] = 1'b0; \
	doodle_left_alpha[40][15] = 1'b0; \
	doodle_left_alpha[40][16] = 1'b0; \
	doodle_left_alpha[40][17] = 1'b0; \
	doodle_left_alpha[40][18] = 1'b0; \
	doodle_left_alpha[40][19] = 1'b0; \
	doodle_left_alpha[40][20] = 1'b0; \
	doodle_left_alpha[40][21] = 1'b0; \
	doodle_left_alpha[40][22] = 1'b0; \
	doodle_left_alpha[40][23] = 1'b0; \
	doodle_left_alpha[40][24] = 1'b0; \
	doodle_left_alpha[40][25] = 1'b0; \
	doodle_left_alpha[40][26] = 1'b0; \
	doodle_left_alpha[40][27] = 1'b0; \
	doodle_left_alpha[40][28] = 1'b0; \
	doodle_left_alpha[40][29] = 1'b0; \
	doodle_left_alpha[40][30] = 1'b0; \
	doodle_left_alpha[40][31] = 1'b0; \
	doodle_left_alpha[40][32] = 1'b0; \
	doodle_left_alpha[40][33] = 1'b0; \
	doodle_left_alpha[40][34] = 1'b0; \
	doodle_left_alpha[40][35] = 1'b0; \
	doodle_left_alpha[40][36] = 1'b0; \
	doodle_left_alpha[40][37] = 1'b0; \
	doodle_left_alpha[40][38] = 1'b0; \
	doodle_left_alpha[40][39] = 1'b0; \
	doodle_left_alpha[40][40] = 1'b0; \
	doodle_left_alpha[40][41] = 1'b0; \
	doodle_left_alpha[40][42] = 1'b0; \
	doodle_left_alpha[40][43] = 1'b0; \
	doodle_left_alpha[40][44] = 1'b0; \
	doodle_left_alpha[40][45] = 1'b0; \
	doodle_left_alpha[40][46] = 1'b0; \
	doodle_left_alpha[40][47] = 1'b0; \
	doodle_left_alpha[40][48] = 1'b0; \
	doodle_left_alpha[40][49] = 1'b0; \
	doodle_left_alpha[40][50] = 1'b0; \
	doodle_left_alpha[40][51] = 1'b0; \
	doodle_left_alpha[40][52] = 1'b0; \
	doodle_left_alpha[40][53] = 1'b0; \
	doodle_left_alpha[40][54] = 1'b0; \
	doodle_left_alpha[40][55] = 1'b0; \
	doodle_left_alpha[40][56] = 1'b0; \
	doodle_left_alpha[40][57] = 1'b0; \
	doodle_left_alpha[40][58] = 1'b0; \
	doodle_left_alpha[40][59] = 1'b0; \
	doodle_left_alpha[40][60] = 1'b0; \
	doodle_left_alpha[40][61] = 1'b0; \
	doodle_left_alpha[40][62] = 1'b0; \
	doodle_left_alpha[40][63] = 1'b0; \
	doodle_left_alpha[40][64] = 1'b0; \
	doodle_left_alpha[40][65] = 1'b1; \
	doodle_left_alpha[40][66] = 1'b1; \
	doodle_left_alpha[40][67] = 1'b1; \
	doodle_left_alpha[40][68] = 1'b1; \
	doodle_left_alpha[40][69] = 1'b1; \
	doodle_left_alpha[40][70] = 1'b1; \
	doodle_left_alpha[40][71] = 1'b1; \
	doodle_left_alpha[40][72] = 1'b1; \
	doodle_left_alpha[40][73] = 1'b1; \
	doodle_left_alpha[40][74] = 1'b1; \
	doodle_left_alpha[40][75] = 1'b1; \
	doodle_left_alpha[40][76] = 1'b1; \
	doodle_left_alpha[40][77] = 1'b1; \
	doodle_left_alpha[40][78] = 1'b1; \
	doodle_left_alpha[40][79] = 1'b1; \
	doodle_left_alpha[41][0] = 1'b1; \
	doodle_left_alpha[41][1] = 1'b1; \
	doodle_left_alpha[41][2] = 1'b1; \
	doodle_left_alpha[41][3] = 1'b1; \
	doodle_left_alpha[41][4] = 1'b0; \
	doodle_left_alpha[41][5] = 1'b0; \
	doodle_left_alpha[41][6] = 1'b0; \
	doodle_left_alpha[41][7] = 1'b0; \
	doodle_left_alpha[41][8] = 1'b0; \
	doodle_left_alpha[41][9] = 1'b0; \
	doodle_left_alpha[41][10] = 1'b0; \
	doodle_left_alpha[41][11] = 1'b0; \
	doodle_left_alpha[41][12] = 1'b0; \
	doodle_left_alpha[41][13] = 1'b0; \
	doodle_left_alpha[41][14] = 1'b0; \
	doodle_left_alpha[41][15] = 1'b0; \
	doodle_left_alpha[41][16] = 1'b0; \
	doodle_left_alpha[41][17] = 1'b0; \
	doodle_left_alpha[41][18] = 1'b0; \
	doodle_left_alpha[41][19] = 1'b0; \
	doodle_left_alpha[41][20] = 1'b0; \
	doodle_left_alpha[41][21] = 1'b0; \
	doodle_left_alpha[41][22] = 1'b0; \
	doodle_left_alpha[41][23] = 1'b0; \
	doodle_left_alpha[41][24] = 1'b0; \
	doodle_left_alpha[41][25] = 1'b0; \
	doodle_left_alpha[41][26] = 1'b0; \
	doodle_left_alpha[41][27] = 1'b0; \
	doodle_left_alpha[41][28] = 1'b0; \
	doodle_left_alpha[41][29] = 1'b0; \
	doodle_left_alpha[41][30] = 1'b0; \
	doodle_left_alpha[41][31] = 1'b0; \
	doodle_left_alpha[41][32] = 1'b0; \
	doodle_left_alpha[41][33] = 1'b0; \
	doodle_left_alpha[41][34] = 1'b0; \
	doodle_left_alpha[41][35] = 1'b0; \
	doodle_left_alpha[41][36] = 1'b0; \
	doodle_left_alpha[41][37] = 1'b0; \
	doodle_left_alpha[41][38] = 1'b0; \
	doodle_left_alpha[41][39] = 1'b0; \
	doodle_left_alpha[41][40] = 1'b0; \
	doodle_left_alpha[41][41] = 1'b0; \
	doodle_left_alpha[41][42] = 1'b0; \
	doodle_left_alpha[41][43] = 1'b0; \
	doodle_left_alpha[41][44] = 1'b0; \
	doodle_left_alpha[41][45] = 1'b0; \
	doodle_left_alpha[41][46] = 1'b0; \
	doodle_left_alpha[41][47] = 1'b0; \
	doodle_left_alpha[41][48] = 1'b0; \
	doodle_left_alpha[41][49] = 1'b0; \
	doodle_left_alpha[41][50] = 1'b0; \
	doodle_left_alpha[41][51] = 1'b0; \
	doodle_left_alpha[41][52] = 1'b0; \
	doodle_left_alpha[41][53] = 1'b0; \
	doodle_left_alpha[41][54] = 1'b0; \
	doodle_left_alpha[41][55] = 1'b0; \
	doodle_left_alpha[41][56] = 1'b0; \
	doodle_left_alpha[41][57] = 1'b0; \
	doodle_left_alpha[41][58] = 1'b0; \
	doodle_left_alpha[41][59] = 1'b0; \
	doodle_left_alpha[41][60] = 1'b0; \
	doodle_left_alpha[41][61] = 1'b0; \
	doodle_left_alpha[41][62] = 1'b0; \
	doodle_left_alpha[41][63] = 1'b0; \
	doodle_left_alpha[41][64] = 1'b0; \
	doodle_left_alpha[41][65] = 1'b1; \
	doodle_left_alpha[41][66] = 1'b1; \
	doodle_left_alpha[41][67] = 1'b1; \
	doodle_left_alpha[41][68] = 1'b1; \
	doodle_left_alpha[41][69] = 1'b1; \
	doodle_left_alpha[41][70] = 1'b1; \
	doodle_left_alpha[41][71] = 1'b1; \
	doodle_left_alpha[41][72] = 1'b1; \
	doodle_left_alpha[41][73] = 1'b1; \
	doodle_left_alpha[41][74] = 1'b1; \
	doodle_left_alpha[41][75] = 1'b1; \
	doodle_left_alpha[41][76] = 1'b1; \
	doodle_left_alpha[41][77] = 1'b1; \
	doodle_left_alpha[41][78] = 1'b1; \
	doodle_left_alpha[41][79] = 1'b1; \
	doodle_left_alpha[42][0] = 1'b1; \
	doodle_left_alpha[42][1] = 1'b1; \
	doodle_left_alpha[42][2] = 1'b1; \
	doodle_left_alpha[42][3] = 1'b1; \
	doodle_left_alpha[42][4] = 1'b0; \
	doodle_left_alpha[42][5] = 1'b0; \
	doodle_left_alpha[42][6] = 1'b0; \
	doodle_left_alpha[42][7] = 1'b0; \
	doodle_left_alpha[42][8] = 1'b0; \
	doodle_left_alpha[42][9] = 1'b0; \
	doodle_left_alpha[42][10] = 1'b0; \
	doodle_left_alpha[42][11] = 1'b0; \
	doodle_left_alpha[42][12] = 1'b0; \
	doodle_left_alpha[42][13] = 1'b0; \
	doodle_left_alpha[42][14] = 1'b0; \
	doodle_left_alpha[42][15] = 1'b0; \
	doodle_left_alpha[42][16] = 1'b0; \
	doodle_left_alpha[42][17] = 1'b0; \
	doodle_left_alpha[42][18] = 1'b0; \
	doodle_left_alpha[42][19] = 1'b0; \
	doodle_left_alpha[42][20] = 1'b0; \
	doodle_left_alpha[42][21] = 1'b0; \
	doodle_left_alpha[42][22] = 1'b0; \
	doodle_left_alpha[42][23] = 1'b0; \
	doodle_left_alpha[42][24] = 1'b0; \
	doodle_left_alpha[42][25] = 1'b0; \
	doodle_left_alpha[42][26] = 1'b0; \
	doodle_left_alpha[42][27] = 1'b0; \
	doodle_left_alpha[42][28] = 1'b0; \
	doodle_left_alpha[42][29] = 1'b0; \
	doodle_left_alpha[42][30] = 1'b0; \
	doodle_left_alpha[42][31] = 1'b0; \
	doodle_left_alpha[42][32] = 1'b0; \
	doodle_left_alpha[42][33] = 1'b0; \
	doodle_left_alpha[42][34] = 1'b0; \
	doodle_left_alpha[42][35] = 1'b0; \
	doodle_left_alpha[42][36] = 1'b0; \
	doodle_left_alpha[42][37] = 1'b0; \
	doodle_left_alpha[42][38] = 1'b0; \
	doodle_left_alpha[42][39] = 1'b0; \
	doodle_left_alpha[42][40] = 1'b0; \
	doodle_left_alpha[42][41] = 1'b0; \
	doodle_left_alpha[42][42] = 1'b0; \
	doodle_left_alpha[42][43] = 1'b0; \
	doodle_left_alpha[42][44] = 1'b0; \
	doodle_left_alpha[42][45] = 1'b0; \
	doodle_left_alpha[42][46] = 1'b0; \
	doodle_left_alpha[42][47] = 1'b0; \
	doodle_left_alpha[42][48] = 1'b0; \
	doodle_left_alpha[42][49] = 1'b0; \
	doodle_left_alpha[42][50] = 1'b0; \
	doodle_left_alpha[42][51] = 1'b0; \
	doodle_left_alpha[42][52] = 1'b0; \
	doodle_left_alpha[42][53] = 1'b0; \
	doodle_left_alpha[42][54] = 1'b0; \
	doodle_left_alpha[42][55] = 1'b0; \
	doodle_left_alpha[42][56] = 1'b0; \
	doodle_left_alpha[42][57] = 1'b0; \
	doodle_left_alpha[42][58] = 1'b0; \
	doodle_left_alpha[42][59] = 1'b0; \
	doodle_left_alpha[42][60] = 1'b0; \
	doodle_left_alpha[42][61] = 1'b0; \
	doodle_left_alpha[42][62] = 1'b0; \
	doodle_left_alpha[42][63] = 1'b0; \
	doodle_left_alpha[42][64] = 1'b0; \
	doodle_left_alpha[42][65] = 1'b1; \
	doodle_left_alpha[42][66] = 1'b1; \
	doodle_left_alpha[42][67] = 1'b1; \
	doodle_left_alpha[42][68] = 1'b1; \
	doodle_left_alpha[42][69] = 1'b1; \
	doodle_left_alpha[42][70] = 1'b1; \
	doodle_left_alpha[42][71] = 1'b1; \
	doodle_left_alpha[42][72] = 1'b1; \
	doodle_left_alpha[42][73] = 1'b1; \
	doodle_left_alpha[42][74] = 1'b1; \
	doodle_left_alpha[42][75] = 1'b1; \
	doodle_left_alpha[42][76] = 1'b1; \
	doodle_left_alpha[42][77] = 1'b1; \
	doodle_left_alpha[42][78] = 1'b1; \
	doodle_left_alpha[42][79] = 1'b1; \
	doodle_left_alpha[43][0] = 1'b1; \
	doodle_left_alpha[43][1] = 1'b1; \
	doodle_left_alpha[43][2] = 1'b1; \
	doodle_left_alpha[43][3] = 1'b1; \
	doodle_left_alpha[43][4] = 1'b0; \
	doodle_left_alpha[43][5] = 1'b0; \
	doodle_left_alpha[43][6] = 1'b0; \
	doodle_left_alpha[43][7] = 1'b0; \
	doodle_left_alpha[43][8] = 1'b0; \
	doodle_left_alpha[43][9] = 1'b0; \
	doodle_left_alpha[43][10] = 1'b0; \
	doodle_left_alpha[43][11] = 1'b0; \
	doodle_left_alpha[43][12] = 1'b0; \
	doodle_left_alpha[43][13] = 1'b0; \
	doodle_left_alpha[43][14] = 1'b0; \
	doodle_left_alpha[43][15] = 1'b0; \
	doodle_left_alpha[43][16] = 1'b0; \
	doodle_left_alpha[43][17] = 1'b0; \
	doodle_left_alpha[43][18] = 1'b0; \
	doodle_left_alpha[43][19] = 1'b0; \
	doodle_left_alpha[43][20] = 1'b0; \
	doodle_left_alpha[43][21] = 1'b0; \
	doodle_left_alpha[43][22] = 1'b0; \
	doodle_left_alpha[43][23] = 1'b0; \
	doodle_left_alpha[43][24] = 1'b0; \
	doodle_left_alpha[43][25] = 1'b0; \
	doodle_left_alpha[43][26] = 1'b0; \
	doodle_left_alpha[43][27] = 1'b0; \
	doodle_left_alpha[43][28] = 1'b0; \
	doodle_left_alpha[43][29] = 1'b0; \
	doodle_left_alpha[43][30] = 1'b0; \
	doodle_left_alpha[43][31] = 1'b0; \
	doodle_left_alpha[43][32] = 1'b0; \
	doodle_left_alpha[43][33] = 1'b0; \
	doodle_left_alpha[43][34] = 1'b0; \
	doodle_left_alpha[43][35] = 1'b0; \
	doodle_left_alpha[43][36] = 1'b0; \
	doodle_left_alpha[43][37] = 1'b0; \
	doodle_left_alpha[43][38] = 1'b0; \
	doodle_left_alpha[43][39] = 1'b0; \
	doodle_left_alpha[43][40] = 1'b0; \
	doodle_left_alpha[43][41] = 1'b0; \
	doodle_left_alpha[43][42] = 1'b0; \
	doodle_left_alpha[43][43] = 1'b0; \
	doodle_left_alpha[43][44] = 1'b0; \
	doodle_left_alpha[43][45] = 1'b0; \
	doodle_left_alpha[43][46] = 1'b0; \
	doodle_left_alpha[43][47] = 1'b0; \
	doodle_left_alpha[43][48] = 1'b0; \
	doodle_left_alpha[43][49] = 1'b0; \
	doodle_left_alpha[43][50] = 1'b0; \
	doodle_left_alpha[43][51] = 1'b0; \
	doodle_left_alpha[43][52] = 1'b0; \
	doodle_left_alpha[43][53] = 1'b0; \
	doodle_left_alpha[43][54] = 1'b0; \
	doodle_left_alpha[43][55] = 1'b0; \
	doodle_left_alpha[43][56] = 1'b0; \
	doodle_left_alpha[43][57] = 1'b0; \
	doodle_left_alpha[43][58] = 1'b0; \
	doodle_left_alpha[43][59] = 1'b0; \
	doodle_left_alpha[43][60] = 1'b0; \
	doodle_left_alpha[43][61] = 1'b0; \
	doodle_left_alpha[43][62] = 1'b0; \
	doodle_left_alpha[43][63] = 1'b0; \
	doodle_left_alpha[43][64] = 1'b0; \
	doodle_left_alpha[43][65] = 1'b1; \
	doodle_left_alpha[43][66] = 1'b1; \
	doodle_left_alpha[43][67] = 1'b1; \
	doodle_left_alpha[43][68] = 1'b1; \
	doodle_left_alpha[43][69] = 1'b1; \
	doodle_left_alpha[43][70] = 1'b1; \
	doodle_left_alpha[43][71] = 1'b1; \
	doodle_left_alpha[43][72] = 1'b1; \
	doodle_left_alpha[43][73] = 1'b1; \
	doodle_left_alpha[43][74] = 1'b1; \
	doodle_left_alpha[43][75] = 1'b1; \
	doodle_left_alpha[43][76] = 1'b1; \
	doodle_left_alpha[43][77] = 1'b1; \
	doodle_left_alpha[43][78] = 1'b1; \
	doodle_left_alpha[43][79] = 1'b1; \
	doodle_left_alpha[44][0] = 1'b1; \
	doodle_left_alpha[44][1] = 1'b1; \
	doodle_left_alpha[44][2] = 1'b1; \
	doodle_left_alpha[44][3] = 1'b1; \
	doodle_left_alpha[44][4] = 1'b0; \
	doodle_left_alpha[44][5] = 1'b0; \
	doodle_left_alpha[44][6] = 1'b0; \
	doodle_left_alpha[44][7] = 1'b0; \
	doodle_left_alpha[44][8] = 1'b0; \
	doodle_left_alpha[44][9] = 1'b0; \
	doodle_left_alpha[44][10] = 1'b0; \
	doodle_left_alpha[44][11] = 1'b0; \
	doodle_left_alpha[44][12] = 1'b0; \
	doodle_left_alpha[44][13] = 1'b0; \
	doodle_left_alpha[44][14] = 1'b0; \
	doodle_left_alpha[44][15] = 1'b0; \
	doodle_left_alpha[44][16] = 1'b0; \
	doodle_left_alpha[44][17] = 1'b0; \
	doodle_left_alpha[44][18] = 1'b0; \
	doodle_left_alpha[44][19] = 1'b0; \
	doodle_left_alpha[44][20] = 1'b0; \
	doodle_left_alpha[44][21] = 1'b0; \
	doodle_left_alpha[44][22] = 1'b0; \
	doodle_left_alpha[44][23] = 1'b0; \
	doodle_left_alpha[44][24] = 1'b0; \
	doodle_left_alpha[44][25] = 1'b0; \
	doodle_left_alpha[44][26] = 1'b0; \
	doodle_left_alpha[44][27] = 1'b0; \
	doodle_left_alpha[44][28] = 1'b0; \
	doodle_left_alpha[44][29] = 1'b0; \
	doodle_left_alpha[44][30] = 1'b0; \
	doodle_left_alpha[44][31] = 1'b0; \
	doodle_left_alpha[44][32] = 1'b0; \
	doodle_left_alpha[44][33] = 1'b0; \
	doodle_left_alpha[44][34] = 1'b0; \
	doodle_left_alpha[44][35] = 1'b0; \
	doodle_left_alpha[44][36] = 1'b0; \
	doodle_left_alpha[44][37] = 1'b0; \
	doodle_left_alpha[44][38] = 1'b0; \
	doodle_left_alpha[44][39] = 1'b0; \
	doodle_left_alpha[44][40] = 1'b0; \
	doodle_left_alpha[44][41] = 1'b0; \
	doodle_left_alpha[44][42] = 1'b0; \
	doodle_left_alpha[44][43] = 1'b0; \
	doodle_left_alpha[44][44] = 1'b0; \
	doodle_left_alpha[44][45] = 1'b0; \
	doodle_left_alpha[44][46] = 1'b0; \
	doodle_left_alpha[44][47] = 1'b0; \
	doodle_left_alpha[44][48] = 1'b0; \
	doodle_left_alpha[44][49] = 1'b0; \
	doodle_left_alpha[44][50] = 1'b0; \
	doodle_left_alpha[44][51] = 1'b0; \
	doodle_left_alpha[44][52] = 1'b0; \
	doodle_left_alpha[44][53] = 1'b0; \
	doodle_left_alpha[44][54] = 1'b0; \
	doodle_left_alpha[44][55] = 1'b0; \
	doodle_left_alpha[44][56] = 1'b0; \
	doodle_left_alpha[44][57] = 1'b0; \
	doodle_left_alpha[44][58] = 1'b0; \
	doodle_left_alpha[44][59] = 1'b0; \
	doodle_left_alpha[44][60] = 1'b0; \
	doodle_left_alpha[44][61] = 1'b0; \
	doodle_left_alpha[44][62] = 1'b0; \
	doodle_left_alpha[44][63] = 1'b0; \
	doodle_left_alpha[44][64] = 1'b0; \
	doodle_left_alpha[44][65] = 1'b1; \
	doodle_left_alpha[44][66] = 1'b1; \
	doodle_left_alpha[44][67] = 1'b1; \
	doodle_left_alpha[44][68] = 1'b1; \
	doodle_left_alpha[44][69] = 1'b1; \
	doodle_left_alpha[44][70] = 1'b1; \
	doodle_left_alpha[44][71] = 1'b1; \
	doodle_left_alpha[44][72] = 1'b1; \
	doodle_left_alpha[44][73] = 1'b1; \
	doodle_left_alpha[44][74] = 1'b1; \
	doodle_left_alpha[44][75] = 1'b1; \
	doodle_left_alpha[44][76] = 1'b1; \
	doodle_left_alpha[44][77] = 1'b1; \
	doodle_left_alpha[44][78] = 1'b1; \
	doodle_left_alpha[44][79] = 1'b1; \
	doodle_left_alpha[45][0] = 1'b1; \
	doodle_left_alpha[45][1] = 1'b1; \
	doodle_left_alpha[45][2] = 1'b1; \
	doodle_left_alpha[45][3] = 1'b1; \
	doodle_left_alpha[45][4] = 1'b0; \
	doodle_left_alpha[45][5] = 1'b0; \
	doodle_left_alpha[45][6] = 1'b0; \
	doodle_left_alpha[45][7] = 1'b0; \
	doodle_left_alpha[45][8] = 1'b0; \
	doodle_left_alpha[45][9] = 1'b0; \
	doodle_left_alpha[45][10] = 1'b0; \
	doodle_left_alpha[45][11] = 1'b0; \
	doodle_left_alpha[45][12] = 1'b0; \
	doodle_left_alpha[45][13] = 1'b0; \
	doodle_left_alpha[45][14] = 1'b0; \
	doodle_left_alpha[45][15] = 1'b0; \
	doodle_left_alpha[45][16] = 1'b0; \
	doodle_left_alpha[45][17] = 1'b0; \
	doodle_left_alpha[45][18] = 1'b0; \
	doodle_left_alpha[45][19] = 1'b0; \
	doodle_left_alpha[45][20] = 1'b0; \
	doodle_left_alpha[45][21] = 1'b0; \
	doodle_left_alpha[45][22] = 1'b0; \
	doodle_left_alpha[45][23] = 1'b0; \
	doodle_left_alpha[45][24] = 1'b0; \
	doodle_left_alpha[45][25] = 1'b0; \
	doodle_left_alpha[45][26] = 1'b0; \
	doodle_left_alpha[45][27] = 1'b0; \
	doodle_left_alpha[45][28] = 1'b0; \
	doodle_left_alpha[45][29] = 1'b0; \
	doodle_left_alpha[45][30] = 1'b0; \
	doodle_left_alpha[45][31] = 1'b0; \
	doodle_left_alpha[45][32] = 1'b0; \
	doodle_left_alpha[45][33] = 1'b0; \
	doodle_left_alpha[45][34] = 1'b0; \
	doodle_left_alpha[45][35] = 1'b0; \
	doodle_left_alpha[45][36] = 1'b0; \
	doodle_left_alpha[45][37] = 1'b0; \
	doodle_left_alpha[45][38] = 1'b0; \
	doodle_left_alpha[45][39] = 1'b0; \
	doodle_left_alpha[45][40] = 1'b0; \
	doodle_left_alpha[45][41] = 1'b0; \
	doodle_left_alpha[45][42] = 1'b0; \
	doodle_left_alpha[45][43] = 1'b0; \
	doodle_left_alpha[45][44] = 1'b0; \
	doodle_left_alpha[45][45] = 1'b0; \
	doodle_left_alpha[45][46] = 1'b0; \
	doodle_left_alpha[45][47] = 1'b0; \
	doodle_left_alpha[45][48] = 1'b0; \
	doodle_left_alpha[45][49] = 1'b0; \
	doodle_left_alpha[45][50] = 1'b0; \
	doodle_left_alpha[45][51] = 1'b0; \
	doodle_left_alpha[45][52] = 1'b0; \
	doodle_left_alpha[45][53] = 1'b0; \
	doodle_left_alpha[45][54] = 1'b0; \
	doodle_left_alpha[45][55] = 1'b0; \
	doodle_left_alpha[45][56] = 1'b0; \
	doodle_left_alpha[45][57] = 1'b0; \
	doodle_left_alpha[45][58] = 1'b0; \
	doodle_left_alpha[45][59] = 1'b0; \
	doodle_left_alpha[45][60] = 1'b0; \
	doodle_left_alpha[45][61] = 1'b0; \
	doodle_left_alpha[45][62] = 1'b0; \
	doodle_left_alpha[45][63] = 1'b0; \
	doodle_left_alpha[45][64] = 1'b0; \
	doodle_left_alpha[45][65] = 1'b1; \
	doodle_left_alpha[45][66] = 1'b1; \
	doodle_left_alpha[45][67] = 1'b1; \
	doodle_left_alpha[45][68] = 1'b1; \
	doodle_left_alpha[45][69] = 1'b1; \
	doodle_left_alpha[45][70] = 1'b1; \
	doodle_left_alpha[45][71] = 1'b1; \
	doodle_left_alpha[45][72] = 1'b1; \
	doodle_left_alpha[45][73] = 1'b1; \
	doodle_left_alpha[45][74] = 1'b1; \
	doodle_left_alpha[45][75] = 1'b1; \
	doodle_left_alpha[45][76] = 1'b1; \
	doodle_left_alpha[45][77] = 1'b1; \
	doodle_left_alpha[45][78] = 1'b1; \
	doodle_left_alpha[45][79] = 1'b1; \
	doodle_left_alpha[46][0] = 1'b1; \
	doodle_left_alpha[46][1] = 1'b1; \
	doodle_left_alpha[46][2] = 1'b1; \
	doodle_left_alpha[46][3] = 1'b1; \
	doodle_left_alpha[46][4] = 1'b1; \
	doodle_left_alpha[46][5] = 1'b1; \
	doodle_left_alpha[46][6] = 1'b1; \
	doodle_left_alpha[46][7] = 1'b1; \
	doodle_left_alpha[46][8] = 1'b1; \
	doodle_left_alpha[46][9] = 1'b1; \
	doodle_left_alpha[46][10] = 1'b1; \
	doodle_left_alpha[46][11] = 1'b1; \
	doodle_left_alpha[46][12] = 1'b1; \
	doodle_left_alpha[46][13] = 1'b1; \
	doodle_left_alpha[46][14] = 1'b1; \
	doodle_left_alpha[46][15] = 1'b1; \
	doodle_left_alpha[46][16] = 1'b1; \
	doodle_left_alpha[46][17] = 1'b1; \
	doodle_left_alpha[46][18] = 1'b1; \
	doodle_left_alpha[46][19] = 1'b1; \
	doodle_left_alpha[46][20] = 1'b1; \
	doodle_left_alpha[46][21] = 1'b1; \
	doodle_left_alpha[46][22] = 1'b1; \
	doodle_left_alpha[46][23] = 1'b0; \
	doodle_left_alpha[46][24] = 1'b0; \
	doodle_left_alpha[46][25] = 1'b0; \
	doodle_left_alpha[46][26] = 1'b0; \
	doodle_left_alpha[46][27] = 1'b0; \
	doodle_left_alpha[46][28] = 1'b0; \
	doodle_left_alpha[46][29] = 1'b0; \
	doodle_left_alpha[46][30] = 1'b0; \
	doodle_left_alpha[46][31] = 1'b0; \
	doodle_left_alpha[46][32] = 1'b0; \
	doodle_left_alpha[46][33] = 1'b0; \
	doodle_left_alpha[46][34] = 1'b0; \
	doodle_left_alpha[46][35] = 1'b0; \
	doodle_left_alpha[46][36] = 1'b0; \
	doodle_left_alpha[46][37] = 1'b0; \
	doodle_left_alpha[46][38] = 1'b0; \
	doodle_left_alpha[46][39] = 1'b0; \
	doodle_left_alpha[46][40] = 1'b0; \
	doodle_left_alpha[46][41] = 1'b0; \
	doodle_left_alpha[46][42] = 1'b0; \
	doodle_left_alpha[46][43] = 1'b0; \
	doodle_left_alpha[46][44] = 1'b0; \
	doodle_left_alpha[46][45] = 1'b0; \
	doodle_left_alpha[46][46] = 1'b0; \
	doodle_left_alpha[46][47] = 1'b0; \
	doodle_left_alpha[46][48] = 1'b0; \
	doodle_left_alpha[46][49] = 1'b0; \
	doodle_left_alpha[46][50] = 1'b0; \
	doodle_left_alpha[46][51] = 1'b0; \
	doodle_left_alpha[46][52] = 1'b0; \
	doodle_left_alpha[46][53] = 1'b0; \
	doodle_left_alpha[46][54] = 1'b0; \
	doodle_left_alpha[46][55] = 1'b0; \
	doodle_left_alpha[46][56] = 1'b0; \
	doodle_left_alpha[46][57] = 1'b0; \
	doodle_left_alpha[46][58] = 1'b0; \
	doodle_left_alpha[46][59] = 1'b0; \
	doodle_left_alpha[46][60] = 1'b0; \
	doodle_left_alpha[46][61] = 1'b0; \
	doodle_left_alpha[46][62] = 1'b0; \
	doodle_left_alpha[46][63] = 1'b0; \
	doodle_left_alpha[46][64] = 1'b0; \
	doodle_left_alpha[46][65] = 1'b1; \
	doodle_left_alpha[46][66] = 1'b1; \
	doodle_left_alpha[46][67] = 1'b1; \
	doodle_left_alpha[46][68] = 1'b1; \
	doodle_left_alpha[46][69] = 1'b1; \
	doodle_left_alpha[46][70] = 1'b1; \
	doodle_left_alpha[46][71] = 1'b1; \
	doodle_left_alpha[46][72] = 1'b1; \
	doodle_left_alpha[46][73] = 1'b1; \
	doodle_left_alpha[46][74] = 1'b1; \
	doodle_left_alpha[46][75] = 1'b1; \
	doodle_left_alpha[46][76] = 1'b1; \
	doodle_left_alpha[46][77] = 1'b1; \
	doodle_left_alpha[46][78] = 1'b1; \
	doodle_left_alpha[46][79] = 1'b1; \
	doodle_left_alpha[47][0] = 1'b1; \
	doodle_left_alpha[47][1] = 1'b1; \
	doodle_left_alpha[47][2] = 1'b1; \
	doodle_left_alpha[47][3] = 1'b1; \
	doodle_left_alpha[47][4] = 1'b1; \
	doodle_left_alpha[47][5] = 1'b1; \
	doodle_left_alpha[47][6] = 1'b1; \
	doodle_left_alpha[47][7] = 1'b1; \
	doodle_left_alpha[47][8] = 1'b1; \
	doodle_left_alpha[47][9] = 1'b1; \
	doodle_left_alpha[47][10] = 1'b1; \
	doodle_left_alpha[47][11] = 1'b1; \
	doodle_left_alpha[47][12] = 1'b1; \
	doodle_left_alpha[47][13] = 1'b1; \
	doodle_left_alpha[47][14] = 1'b1; \
	doodle_left_alpha[47][15] = 1'b1; \
	doodle_left_alpha[47][16] = 1'b1; \
	doodle_left_alpha[47][17] = 1'b1; \
	doodle_left_alpha[47][18] = 1'b1; \
	doodle_left_alpha[47][19] = 1'b1; \
	doodle_left_alpha[47][20] = 1'b1; \
	doodle_left_alpha[47][21] = 1'b1; \
	doodle_left_alpha[47][22] = 1'b1; \
	doodle_left_alpha[47][23] = 1'b0; \
	doodle_left_alpha[47][24] = 1'b0; \
	doodle_left_alpha[47][25] = 1'b0; \
	doodle_left_alpha[47][26] = 1'b0; \
	doodle_left_alpha[47][27] = 1'b0; \
	doodle_left_alpha[47][28] = 1'b0; \
	doodle_left_alpha[47][29] = 1'b0; \
	doodle_left_alpha[47][30] = 1'b0; \
	doodle_left_alpha[47][31] = 1'b0; \
	doodle_left_alpha[47][32] = 1'b0; \
	doodle_left_alpha[47][33] = 1'b0; \
	doodle_left_alpha[47][34] = 1'b0; \
	doodle_left_alpha[47][35] = 1'b0; \
	doodle_left_alpha[47][36] = 1'b0; \
	doodle_left_alpha[47][37] = 1'b0; \
	doodle_left_alpha[47][38] = 1'b0; \
	doodle_left_alpha[47][39] = 1'b0; \
	doodle_left_alpha[47][40] = 1'b0; \
	doodle_left_alpha[47][41] = 1'b0; \
	doodle_left_alpha[47][42] = 1'b0; \
	doodle_left_alpha[47][43] = 1'b0; \
	doodle_left_alpha[47][44] = 1'b0; \
	doodle_left_alpha[47][45] = 1'b0; \
	doodle_left_alpha[47][46] = 1'b0; \
	doodle_left_alpha[47][47] = 1'b0; \
	doodle_left_alpha[47][48] = 1'b0; \
	doodle_left_alpha[47][49] = 1'b0; \
	doodle_left_alpha[47][50] = 1'b0; \
	doodle_left_alpha[47][51] = 1'b0; \
	doodle_left_alpha[47][52] = 1'b0; \
	doodle_left_alpha[47][53] = 1'b0; \
	doodle_left_alpha[47][54] = 1'b0; \
	doodle_left_alpha[47][55] = 1'b0; \
	doodle_left_alpha[47][56] = 1'b0; \
	doodle_left_alpha[47][57] = 1'b0; \
	doodle_left_alpha[47][58] = 1'b0; \
	doodle_left_alpha[47][59] = 1'b0; \
	doodle_left_alpha[47][60] = 1'b0; \
	doodle_left_alpha[47][61] = 1'b0; \
	doodle_left_alpha[47][62] = 1'b0; \
	doodle_left_alpha[47][63] = 1'b0; \
	doodle_left_alpha[47][64] = 1'b0; \
	doodle_left_alpha[47][65] = 1'b1; \
	doodle_left_alpha[47][66] = 1'b1; \
	doodle_left_alpha[47][67] = 1'b1; \
	doodle_left_alpha[47][68] = 1'b1; \
	doodle_left_alpha[47][69] = 1'b1; \
	doodle_left_alpha[47][70] = 1'b1; \
	doodle_left_alpha[47][71] = 1'b1; \
	doodle_left_alpha[47][72] = 1'b1; \
	doodle_left_alpha[47][73] = 1'b1; \
	doodle_left_alpha[47][74] = 1'b1; \
	doodle_left_alpha[47][75] = 1'b1; \
	doodle_left_alpha[47][76] = 1'b1; \
	doodle_left_alpha[47][77] = 1'b1; \
	doodle_left_alpha[47][78] = 1'b1; \
	doodle_left_alpha[47][79] = 1'b1; \
	doodle_left_alpha[48][0] = 1'b1; \
	doodle_left_alpha[48][1] = 1'b1; \
	doodle_left_alpha[48][2] = 1'b1; \
	doodle_left_alpha[48][3] = 1'b1; \
	doodle_left_alpha[48][4] = 1'b1; \
	doodle_left_alpha[48][5] = 1'b1; \
	doodle_left_alpha[48][6] = 1'b1; \
	doodle_left_alpha[48][7] = 1'b1; \
	doodle_left_alpha[48][8] = 1'b1; \
	doodle_left_alpha[48][9] = 1'b1; \
	doodle_left_alpha[48][10] = 1'b1; \
	doodle_left_alpha[48][11] = 1'b1; \
	doodle_left_alpha[48][12] = 1'b1; \
	doodle_left_alpha[48][13] = 1'b1; \
	doodle_left_alpha[48][14] = 1'b1; \
	doodle_left_alpha[48][15] = 1'b1; \
	doodle_left_alpha[48][16] = 1'b1; \
	doodle_left_alpha[48][17] = 1'b1; \
	doodle_left_alpha[48][18] = 1'b1; \
	doodle_left_alpha[48][19] = 1'b1; \
	doodle_left_alpha[48][20] = 1'b1; \
	doodle_left_alpha[48][21] = 1'b1; \
	doodle_left_alpha[48][22] = 1'b1; \
	doodle_left_alpha[48][23] = 1'b0; \
	doodle_left_alpha[48][24] = 1'b0; \
	doodle_left_alpha[48][25] = 1'b0; \
	doodle_left_alpha[48][26] = 1'b0; \
	doodle_left_alpha[48][27] = 1'b0; \
	doodle_left_alpha[48][28] = 1'b0; \
	doodle_left_alpha[48][29] = 1'b0; \
	doodle_left_alpha[48][30] = 1'b0; \
	doodle_left_alpha[48][31] = 1'b0; \
	doodle_left_alpha[48][32] = 1'b0; \
	doodle_left_alpha[48][33] = 1'b0; \
	doodle_left_alpha[48][34] = 1'b0; \
	doodle_left_alpha[48][35] = 1'b0; \
	doodle_left_alpha[48][36] = 1'b0; \
	doodle_left_alpha[48][37] = 1'b0; \
	doodle_left_alpha[48][38] = 1'b0; \
	doodle_left_alpha[48][39] = 1'b0; \
	doodle_left_alpha[48][40] = 1'b0; \
	doodle_left_alpha[48][41] = 1'b0; \
	doodle_left_alpha[48][42] = 1'b0; \
	doodle_left_alpha[48][43] = 1'b0; \
	doodle_left_alpha[48][44] = 1'b0; \
	doodle_left_alpha[48][45] = 1'b0; \
	doodle_left_alpha[48][46] = 1'b0; \
	doodle_left_alpha[48][47] = 1'b0; \
	doodle_left_alpha[48][48] = 1'b0; \
	doodle_left_alpha[48][49] = 1'b0; \
	doodle_left_alpha[48][50] = 1'b0; \
	doodle_left_alpha[48][51] = 1'b0; \
	doodle_left_alpha[48][52] = 1'b0; \
	doodle_left_alpha[48][53] = 1'b0; \
	doodle_left_alpha[48][54] = 1'b0; \
	doodle_left_alpha[48][55] = 1'b0; \
	doodle_left_alpha[48][56] = 1'b0; \
	doodle_left_alpha[48][57] = 1'b0; \
	doodle_left_alpha[48][58] = 1'b0; \
	doodle_left_alpha[48][59] = 1'b0; \
	doodle_left_alpha[48][60] = 1'b0; \
	doodle_left_alpha[48][61] = 1'b0; \
	doodle_left_alpha[48][62] = 1'b0; \
	doodle_left_alpha[48][63] = 1'b0; \
	doodle_left_alpha[48][64] = 1'b0; \
	doodle_left_alpha[48][65] = 1'b1; \
	doodle_left_alpha[48][66] = 1'b1; \
	doodle_left_alpha[48][67] = 1'b1; \
	doodle_left_alpha[48][68] = 1'b1; \
	doodle_left_alpha[48][69] = 1'b1; \
	doodle_left_alpha[48][70] = 1'b1; \
	doodle_left_alpha[48][71] = 1'b1; \
	doodle_left_alpha[48][72] = 1'b1; \
	doodle_left_alpha[48][73] = 1'b1; \
	doodle_left_alpha[48][74] = 1'b1; \
	doodle_left_alpha[48][75] = 1'b1; \
	doodle_left_alpha[48][76] = 1'b1; \
	doodle_left_alpha[48][77] = 1'b1; \
	doodle_left_alpha[48][78] = 1'b1; \
	doodle_left_alpha[48][79] = 1'b1; \
	doodle_left_alpha[49][0] = 1'b1; \
	doodle_left_alpha[49][1] = 1'b1; \
	doodle_left_alpha[49][2] = 1'b1; \
	doodle_left_alpha[49][3] = 1'b1; \
	doodle_left_alpha[49][4] = 1'b1; \
	doodle_left_alpha[49][5] = 1'b1; \
	doodle_left_alpha[49][6] = 1'b1; \
	doodle_left_alpha[49][7] = 1'b1; \
	doodle_left_alpha[49][8] = 1'b1; \
	doodle_left_alpha[49][9] = 1'b1; \
	doodle_left_alpha[49][10] = 1'b1; \
	doodle_left_alpha[49][11] = 1'b1; \
	doodle_left_alpha[49][12] = 1'b1; \
	doodle_left_alpha[49][13] = 1'b1; \
	doodle_left_alpha[49][14] = 1'b1; \
	doodle_left_alpha[49][15] = 1'b1; \
	doodle_left_alpha[49][16] = 1'b1; \
	doodle_left_alpha[49][17] = 1'b1; \
	doodle_left_alpha[49][18] = 1'b1; \
	doodle_left_alpha[49][19] = 1'b1; \
	doodle_left_alpha[49][20] = 1'b1; \
	doodle_left_alpha[49][21] = 1'b1; \
	doodle_left_alpha[49][22] = 1'b1; \
	doodle_left_alpha[49][23] = 1'b0; \
	doodle_left_alpha[49][24] = 1'b0; \
	doodle_left_alpha[49][25] = 1'b0; \
	doodle_left_alpha[49][26] = 1'b0; \
	doodle_left_alpha[49][27] = 1'b0; \
	doodle_left_alpha[49][28] = 1'b0; \
	doodle_left_alpha[49][29] = 1'b0; \
	doodle_left_alpha[49][30] = 1'b0; \
	doodle_left_alpha[49][31] = 1'b0; \
	doodle_left_alpha[49][32] = 1'b0; \
	doodle_left_alpha[49][33] = 1'b0; \
	doodle_left_alpha[49][34] = 1'b0; \
	doodle_left_alpha[49][35] = 1'b0; \
	doodle_left_alpha[49][36] = 1'b0; \
	doodle_left_alpha[49][37] = 1'b0; \
	doodle_left_alpha[49][38] = 1'b0; \
	doodle_left_alpha[49][39] = 1'b0; \
	doodle_left_alpha[49][40] = 1'b0; \
	doodle_left_alpha[49][41] = 1'b0; \
	doodle_left_alpha[49][42] = 1'b0; \
	doodle_left_alpha[49][43] = 1'b0; \
	doodle_left_alpha[49][44] = 1'b0; \
	doodle_left_alpha[49][45] = 1'b0; \
	doodle_left_alpha[49][46] = 1'b0; \
	doodle_left_alpha[49][47] = 1'b0; \
	doodle_left_alpha[49][48] = 1'b0; \
	doodle_left_alpha[49][49] = 1'b0; \
	doodle_left_alpha[49][50] = 1'b0; \
	doodle_left_alpha[49][51] = 1'b0; \
	doodle_left_alpha[49][52] = 1'b0; \
	doodle_left_alpha[49][53] = 1'b0; \
	doodle_left_alpha[49][54] = 1'b0; \
	doodle_left_alpha[49][55] = 1'b0; \
	doodle_left_alpha[49][56] = 1'b0; \
	doodle_left_alpha[49][57] = 1'b0; \
	doodle_left_alpha[49][58] = 1'b0; \
	doodle_left_alpha[49][59] = 1'b0; \
	doodle_left_alpha[49][60] = 1'b0; \
	doodle_left_alpha[49][61] = 1'b0; \
	doodle_left_alpha[49][62] = 1'b0; \
	doodle_left_alpha[49][63] = 1'b0; \
	doodle_left_alpha[49][64] = 1'b0; \
	doodle_left_alpha[49][65] = 1'b1; \
	doodle_left_alpha[49][66] = 1'b1; \
	doodle_left_alpha[49][67] = 1'b1; \
	doodle_left_alpha[49][68] = 1'b1; \
	doodle_left_alpha[49][69] = 1'b1; \
	doodle_left_alpha[49][70] = 1'b1; \
	doodle_left_alpha[49][71] = 1'b1; \
	doodle_left_alpha[49][72] = 1'b1; \
	doodle_left_alpha[49][73] = 1'b1; \
	doodle_left_alpha[49][74] = 1'b1; \
	doodle_left_alpha[49][75] = 1'b1; \
	doodle_left_alpha[49][76] = 1'b1; \
	doodle_left_alpha[49][77] = 1'b1; \
	doodle_left_alpha[49][78] = 1'b1; \
	doodle_left_alpha[49][79] = 1'b1; \
	doodle_left_alpha[50][0] = 1'b1; \
	doodle_left_alpha[50][1] = 1'b1; \
	doodle_left_alpha[50][2] = 1'b1; \
	doodle_left_alpha[50][3] = 1'b1; \
	doodle_left_alpha[50][4] = 1'b1; \
	doodle_left_alpha[50][5] = 1'b1; \
	doodle_left_alpha[50][6] = 1'b1; \
	doodle_left_alpha[50][7] = 1'b1; \
	doodle_left_alpha[50][8] = 1'b1; \
	doodle_left_alpha[50][9] = 1'b1; \
	doodle_left_alpha[50][10] = 1'b1; \
	doodle_left_alpha[50][11] = 1'b1; \
	doodle_left_alpha[50][12] = 1'b1; \
	doodle_left_alpha[50][13] = 1'b1; \
	doodle_left_alpha[50][14] = 1'b1; \
	doodle_left_alpha[50][15] = 1'b1; \
	doodle_left_alpha[50][16] = 1'b1; \
	doodle_left_alpha[50][17] = 1'b1; \
	doodle_left_alpha[50][18] = 1'b1; \
	doodle_left_alpha[50][19] = 1'b1; \
	doodle_left_alpha[50][20] = 1'b1; \
	doodle_left_alpha[50][21] = 1'b1; \
	doodle_left_alpha[50][22] = 1'b1; \
	doodle_left_alpha[50][23] = 1'b0; \
	doodle_left_alpha[50][24] = 1'b0; \
	doodle_left_alpha[50][25] = 1'b0; \
	doodle_left_alpha[50][26] = 1'b0; \
	doodle_left_alpha[50][27] = 1'b0; \
	doodle_left_alpha[50][28] = 1'b0; \
	doodle_left_alpha[50][29] = 1'b0; \
	doodle_left_alpha[50][30] = 1'b0; \
	doodle_left_alpha[50][31] = 1'b0; \
	doodle_left_alpha[50][32] = 1'b0; \
	doodle_left_alpha[50][33] = 1'b0; \
	doodle_left_alpha[50][34] = 1'b0; \
	doodle_left_alpha[50][35] = 1'b0; \
	doodle_left_alpha[50][36] = 1'b0; \
	doodle_left_alpha[50][37] = 1'b0; \
	doodle_left_alpha[50][38] = 1'b0; \
	doodle_left_alpha[50][39] = 1'b0; \
	doodle_left_alpha[50][40] = 1'b0; \
	doodle_left_alpha[50][41] = 1'b0; \
	doodle_left_alpha[50][42] = 1'b0; \
	doodle_left_alpha[50][43] = 1'b0; \
	doodle_left_alpha[50][44] = 1'b0; \
	doodle_left_alpha[50][45] = 1'b0; \
	doodle_left_alpha[50][46] = 1'b0; \
	doodle_left_alpha[50][47] = 1'b0; \
	doodle_left_alpha[50][48] = 1'b0; \
	doodle_left_alpha[50][49] = 1'b0; \
	doodle_left_alpha[50][50] = 1'b0; \
	doodle_left_alpha[50][51] = 1'b0; \
	doodle_left_alpha[50][52] = 1'b0; \
	doodle_left_alpha[50][53] = 1'b0; \
	doodle_left_alpha[50][54] = 1'b0; \
	doodle_left_alpha[50][55] = 1'b0; \
	doodle_left_alpha[50][56] = 1'b0; \
	doodle_left_alpha[50][57] = 1'b0; \
	doodle_left_alpha[50][58] = 1'b0; \
	doodle_left_alpha[50][59] = 1'b0; \
	doodle_left_alpha[50][60] = 1'b0; \
	doodle_left_alpha[50][61] = 1'b0; \
	doodle_left_alpha[50][62] = 1'b0; \
	doodle_left_alpha[50][63] = 1'b0; \
	doodle_left_alpha[50][64] = 1'b0; \
	doodle_left_alpha[50][65] = 1'b1; \
	doodle_left_alpha[50][66] = 1'b1; \
	doodle_left_alpha[50][67] = 1'b1; \
	doodle_left_alpha[50][68] = 1'b1; \
	doodle_left_alpha[50][69] = 1'b1; \
	doodle_left_alpha[50][70] = 1'b1; \
	doodle_left_alpha[50][71] = 1'b1; \
	doodle_left_alpha[50][72] = 1'b1; \
	doodle_left_alpha[50][73] = 1'b1; \
	doodle_left_alpha[50][74] = 1'b1; \
	doodle_left_alpha[50][75] = 1'b1; \
	doodle_left_alpha[50][76] = 1'b1; \
	doodle_left_alpha[50][77] = 1'b1; \
	doodle_left_alpha[50][78] = 1'b1; \
	doodle_left_alpha[50][79] = 1'b1; \
	doodle_left_alpha[51][0] = 1'b1; \
	doodle_left_alpha[51][1] = 1'b1; \
	doodle_left_alpha[51][2] = 1'b1; \
	doodle_left_alpha[51][3] = 1'b1; \
	doodle_left_alpha[51][4] = 1'b1; \
	doodle_left_alpha[51][5] = 1'b1; \
	doodle_left_alpha[51][6] = 1'b1; \
	doodle_left_alpha[51][7] = 1'b1; \
	doodle_left_alpha[51][8] = 1'b1; \
	doodle_left_alpha[51][9] = 1'b1; \
	doodle_left_alpha[51][10] = 1'b1; \
	doodle_left_alpha[51][11] = 1'b1; \
	doodle_left_alpha[51][12] = 1'b1; \
	doodle_left_alpha[51][13] = 1'b1; \
	doodle_left_alpha[51][14] = 1'b1; \
	doodle_left_alpha[51][15] = 1'b1; \
	doodle_left_alpha[51][16] = 1'b1; \
	doodle_left_alpha[51][17] = 1'b1; \
	doodle_left_alpha[51][18] = 1'b1; \
	doodle_left_alpha[51][19] = 1'b1; \
	doodle_left_alpha[51][20] = 1'b1; \
	doodle_left_alpha[51][21] = 1'b1; \
	doodle_left_alpha[51][22] = 1'b1; \
	doodle_left_alpha[51][23] = 1'b0; \
	doodle_left_alpha[51][24] = 1'b0; \
	doodle_left_alpha[51][25] = 1'b0; \
	doodle_left_alpha[51][26] = 1'b0; \
	doodle_left_alpha[51][27] = 1'b0; \
	doodle_left_alpha[51][28] = 1'b0; \
	doodle_left_alpha[51][29] = 1'b0; \
	doodle_left_alpha[51][30] = 1'b0; \
	doodle_left_alpha[51][31] = 1'b0; \
	doodle_left_alpha[51][32] = 1'b0; \
	doodle_left_alpha[51][33] = 1'b0; \
	doodle_left_alpha[51][34] = 1'b0; \
	doodle_left_alpha[51][35] = 1'b0; \
	doodle_left_alpha[51][36] = 1'b0; \
	doodle_left_alpha[51][37] = 1'b0; \
	doodle_left_alpha[51][38] = 1'b0; \
	doodle_left_alpha[51][39] = 1'b0; \
	doodle_left_alpha[51][40] = 1'b0; \
	doodle_left_alpha[51][41] = 1'b0; \
	doodle_left_alpha[51][42] = 1'b0; \
	doodle_left_alpha[51][43] = 1'b0; \
	doodle_left_alpha[51][44] = 1'b0; \
	doodle_left_alpha[51][45] = 1'b0; \
	doodle_left_alpha[51][46] = 1'b0; \
	doodle_left_alpha[51][47] = 1'b0; \
	doodle_left_alpha[51][48] = 1'b0; \
	doodle_left_alpha[51][49] = 1'b0; \
	doodle_left_alpha[51][50] = 1'b0; \
	doodle_left_alpha[51][51] = 1'b0; \
	doodle_left_alpha[51][52] = 1'b0; \
	doodle_left_alpha[51][53] = 1'b0; \
	doodle_left_alpha[51][54] = 1'b0; \
	doodle_left_alpha[51][55] = 1'b0; \
	doodle_left_alpha[51][56] = 1'b0; \
	doodle_left_alpha[51][57] = 1'b0; \
	doodle_left_alpha[51][58] = 1'b0; \
	doodle_left_alpha[51][59] = 1'b0; \
	doodle_left_alpha[51][60] = 1'b0; \
	doodle_left_alpha[51][61] = 1'b0; \
	doodle_left_alpha[51][62] = 1'b0; \
	doodle_left_alpha[51][63] = 1'b0; \
	doodle_left_alpha[51][64] = 1'b0; \
	doodle_left_alpha[51][65] = 1'b1; \
	doodle_left_alpha[51][66] = 1'b1; \
	doodle_left_alpha[51][67] = 1'b1; \
	doodle_left_alpha[51][68] = 1'b1; \
	doodle_left_alpha[51][69] = 1'b1; \
	doodle_left_alpha[51][70] = 1'b1; \
	doodle_left_alpha[51][71] = 1'b1; \
	doodle_left_alpha[51][72] = 1'b1; \
	doodle_left_alpha[51][73] = 1'b1; \
	doodle_left_alpha[51][74] = 1'b1; \
	doodle_left_alpha[51][75] = 1'b1; \
	doodle_left_alpha[51][76] = 1'b1; \
	doodle_left_alpha[51][77] = 1'b1; \
	doodle_left_alpha[51][78] = 1'b1; \
	doodle_left_alpha[51][79] = 1'b1; \
	doodle_left_alpha[52][0] = 1'b1; \
	doodle_left_alpha[52][1] = 1'b1; \
	doodle_left_alpha[52][2] = 1'b1; \
	doodle_left_alpha[52][3] = 1'b1; \
	doodle_left_alpha[52][4] = 1'b1; \
	doodle_left_alpha[52][5] = 1'b1; \
	doodle_left_alpha[52][6] = 1'b1; \
	doodle_left_alpha[52][7] = 1'b1; \
	doodle_left_alpha[52][8] = 1'b1; \
	doodle_left_alpha[52][9] = 1'b1; \
	doodle_left_alpha[52][10] = 1'b1; \
	doodle_left_alpha[52][11] = 1'b1; \
	doodle_left_alpha[52][12] = 1'b1; \
	doodle_left_alpha[52][13] = 1'b1; \
	doodle_left_alpha[52][14] = 1'b1; \
	doodle_left_alpha[52][15] = 1'b1; \
	doodle_left_alpha[52][16] = 1'b1; \
	doodle_left_alpha[52][17] = 1'b1; \
	doodle_left_alpha[52][18] = 1'b1; \
	doodle_left_alpha[52][19] = 1'b1; \
	doodle_left_alpha[52][20] = 1'b1; \
	doodle_left_alpha[52][21] = 1'b1; \
	doodle_left_alpha[52][22] = 1'b1; \
	doodle_left_alpha[52][23] = 1'b0; \
	doodle_left_alpha[52][24] = 1'b0; \
	doodle_left_alpha[52][25] = 1'b0; \
	doodle_left_alpha[52][26] = 1'b0; \
	doodle_left_alpha[52][27] = 1'b0; \
	doodle_left_alpha[52][28] = 1'b0; \
	doodle_left_alpha[52][29] = 1'b0; \
	doodle_left_alpha[52][30] = 1'b0; \
	doodle_left_alpha[52][31] = 1'b0; \
	doodle_left_alpha[52][32] = 1'b0; \
	doodle_left_alpha[52][33] = 1'b0; \
	doodle_left_alpha[52][34] = 1'b0; \
	doodle_left_alpha[52][35] = 1'b0; \
	doodle_left_alpha[52][36] = 1'b0; \
	doodle_left_alpha[52][37] = 1'b0; \
	doodle_left_alpha[52][38] = 1'b0; \
	doodle_left_alpha[52][39] = 1'b0; \
	doodle_left_alpha[52][40] = 1'b0; \
	doodle_left_alpha[52][41] = 1'b0; \
	doodle_left_alpha[52][42] = 1'b0; \
	doodle_left_alpha[52][43] = 1'b0; \
	doodle_left_alpha[52][44] = 1'b0; \
	doodle_left_alpha[52][45] = 1'b0; \
	doodle_left_alpha[52][46] = 1'b0; \
	doodle_left_alpha[52][47] = 1'b0; \
	doodle_left_alpha[52][48] = 1'b0; \
	doodle_left_alpha[52][49] = 1'b0; \
	doodle_left_alpha[52][50] = 1'b0; \
	doodle_left_alpha[52][51] = 1'b0; \
	doodle_left_alpha[52][52] = 1'b0; \
	doodle_left_alpha[52][53] = 1'b0; \
	doodle_left_alpha[52][54] = 1'b0; \
	doodle_left_alpha[52][55] = 1'b0; \
	doodle_left_alpha[52][56] = 1'b0; \
	doodle_left_alpha[52][57] = 1'b0; \
	doodle_left_alpha[52][58] = 1'b0; \
	doodle_left_alpha[52][59] = 1'b0; \
	doodle_left_alpha[52][60] = 1'b0; \
	doodle_left_alpha[52][61] = 1'b0; \
	doodle_left_alpha[52][62] = 1'b0; \
	doodle_left_alpha[52][63] = 1'b0; \
	doodle_left_alpha[52][64] = 1'b0; \
	doodle_left_alpha[52][65] = 1'b1; \
	doodle_left_alpha[52][66] = 1'b1; \
	doodle_left_alpha[52][67] = 1'b1; \
	doodle_left_alpha[52][68] = 1'b1; \
	doodle_left_alpha[52][69] = 1'b1; \
	doodle_left_alpha[52][70] = 1'b1; \
	doodle_left_alpha[52][71] = 1'b1; \
	doodle_left_alpha[52][72] = 1'b1; \
	doodle_left_alpha[52][73] = 1'b1; \
	doodle_left_alpha[52][74] = 1'b1; \
	doodle_left_alpha[52][75] = 1'b1; \
	doodle_left_alpha[52][76] = 1'b1; \
	doodle_left_alpha[52][77] = 1'b1; \
	doodle_left_alpha[52][78] = 1'b1; \
	doodle_left_alpha[52][79] = 1'b1; \
	doodle_left_alpha[53][0] = 1'b1; \
	doodle_left_alpha[53][1] = 1'b1; \
	doodle_left_alpha[53][2] = 1'b1; \
	doodle_left_alpha[53][3] = 1'b1; \
	doodle_left_alpha[53][4] = 1'b1; \
	doodle_left_alpha[53][5] = 1'b1; \
	doodle_left_alpha[53][6] = 1'b1; \
	doodle_left_alpha[53][7] = 1'b1; \
	doodle_left_alpha[53][8] = 1'b1; \
	doodle_left_alpha[53][9] = 1'b1; \
	doodle_left_alpha[53][10] = 1'b1; \
	doodle_left_alpha[53][11] = 1'b1; \
	doodle_left_alpha[53][12] = 1'b1; \
	doodle_left_alpha[53][13] = 1'b1; \
	doodle_left_alpha[53][14] = 1'b1; \
	doodle_left_alpha[53][15] = 1'b1; \
	doodle_left_alpha[53][16] = 1'b1; \
	doodle_left_alpha[53][17] = 1'b1; \
	doodle_left_alpha[53][18] = 1'b1; \
	doodle_left_alpha[53][19] = 1'b1; \
	doodle_left_alpha[53][20] = 1'b1; \
	doodle_left_alpha[53][21] = 1'b1; \
	doodle_left_alpha[53][22] = 1'b1; \
	doodle_left_alpha[53][23] = 1'b0; \
	doodle_left_alpha[53][24] = 1'b0; \
	doodle_left_alpha[53][25] = 1'b0; \
	doodle_left_alpha[53][26] = 1'b0; \
	doodle_left_alpha[53][27] = 1'b0; \
	doodle_left_alpha[53][28] = 1'b0; \
	doodle_left_alpha[53][29] = 1'b0; \
	doodle_left_alpha[53][30] = 1'b0; \
	doodle_left_alpha[53][31] = 1'b0; \
	doodle_left_alpha[53][32] = 1'b0; \
	doodle_left_alpha[53][33] = 1'b0; \
	doodle_left_alpha[53][34] = 1'b0; \
	doodle_left_alpha[53][35] = 1'b0; \
	doodle_left_alpha[53][36] = 1'b0; \
	doodle_left_alpha[53][37] = 1'b0; \
	doodle_left_alpha[53][38] = 1'b0; \
	doodle_left_alpha[53][39] = 1'b0; \
	doodle_left_alpha[53][40] = 1'b0; \
	doodle_left_alpha[53][41] = 1'b0; \
	doodle_left_alpha[53][42] = 1'b0; \
	doodle_left_alpha[53][43] = 1'b0; \
	doodle_left_alpha[53][44] = 1'b0; \
	doodle_left_alpha[53][45] = 1'b0; \
	doodle_left_alpha[53][46] = 1'b0; \
	doodle_left_alpha[53][47] = 1'b0; \
	doodle_left_alpha[53][48] = 1'b0; \
	doodle_left_alpha[53][49] = 1'b0; \
	doodle_left_alpha[53][50] = 1'b0; \
	doodle_left_alpha[53][51] = 1'b0; \
	doodle_left_alpha[53][52] = 1'b0; \
	doodle_left_alpha[53][53] = 1'b0; \
	doodle_left_alpha[53][54] = 1'b0; \
	doodle_left_alpha[53][55] = 1'b0; \
	doodle_left_alpha[53][56] = 1'b0; \
	doodle_left_alpha[53][57] = 1'b0; \
	doodle_left_alpha[53][58] = 1'b0; \
	doodle_left_alpha[53][59] = 1'b0; \
	doodle_left_alpha[53][60] = 1'b0; \
	doodle_left_alpha[53][61] = 1'b0; \
	doodle_left_alpha[53][62] = 1'b0; \
	doodle_left_alpha[53][63] = 1'b0; \
	doodle_left_alpha[53][64] = 1'b0; \
	doodle_left_alpha[53][65] = 1'b1; \
	doodle_left_alpha[53][66] = 1'b1; \
	doodle_left_alpha[53][67] = 1'b1; \
	doodle_left_alpha[53][68] = 1'b1; \
	doodle_left_alpha[53][69] = 1'b1; \
	doodle_left_alpha[53][70] = 1'b1; \
	doodle_left_alpha[53][71] = 1'b1; \
	doodle_left_alpha[53][72] = 1'b1; \
	doodle_left_alpha[53][73] = 1'b1; \
	doodle_left_alpha[53][74] = 1'b1; \
	doodle_left_alpha[53][75] = 1'b1; \
	doodle_left_alpha[53][76] = 1'b1; \
	doodle_left_alpha[53][77] = 1'b1; \
	doodle_left_alpha[53][78] = 1'b1; \
	doodle_left_alpha[53][79] = 1'b1; \
	doodle_left_alpha[54][0] = 1'b1; \
	doodle_left_alpha[54][1] = 1'b1; \
	doodle_left_alpha[54][2] = 1'b1; \
	doodle_left_alpha[54][3] = 1'b1; \
	doodle_left_alpha[54][4] = 1'b1; \
	doodle_left_alpha[54][5] = 1'b1; \
	doodle_left_alpha[54][6] = 1'b1; \
	doodle_left_alpha[54][7] = 1'b1; \
	doodle_left_alpha[54][8] = 1'b1; \
	doodle_left_alpha[54][9] = 1'b1; \
	doodle_left_alpha[54][10] = 1'b1; \
	doodle_left_alpha[54][11] = 1'b1; \
	doodle_left_alpha[54][12] = 1'b1; \
	doodle_left_alpha[54][13] = 1'b1; \
	doodle_left_alpha[54][14] = 1'b1; \
	doodle_left_alpha[54][15] = 1'b1; \
	doodle_left_alpha[54][16] = 1'b1; \
	doodle_left_alpha[54][17] = 1'b1; \
	doodle_left_alpha[54][18] = 1'b1; \
	doodle_left_alpha[54][19] = 1'b1; \
	doodle_left_alpha[54][20] = 1'b1; \
	doodle_left_alpha[54][21] = 1'b1; \
	doodle_left_alpha[54][22] = 1'b1; \
	doodle_left_alpha[54][23] = 1'b0; \
	doodle_left_alpha[54][24] = 1'b0; \
	doodle_left_alpha[54][25] = 1'b0; \
	doodle_left_alpha[54][26] = 1'b0; \
	doodle_left_alpha[54][27] = 1'b0; \
	doodle_left_alpha[54][28] = 1'b0; \
	doodle_left_alpha[54][29] = 1'b0; \
	doodle_left_alpha[54][30] = 1'b0; \
	doodle_left_alpha[54][31] = 1'b0; \
	doodle_left_alpha[54][32] = 1'b0; \
	doodle_left_alpha[54][33] = 1'b0; \
	doodle_left_alpha[54][34] = 1'b0; \
	doodle_left_alpha[54][35] = 1'b0; \
	doodle_left_alpha[54][36] = 1'b0; \
	doodle_left_alpha[54][37] = 1'b0; \
	doodle_left_alpha[54][38] = 1'b0; \
	doodle_left_alpha[54][39] = 1'b0; \
	doodle_left_alpha[54][40] = 1'b0; \
	doodle_left_alpha[54][41] = 1'b0; \
	doodle_left_alpha[54][42] = 1'b0; \
	doodle_left_alpha[54][43] = 1'b0; \
	doodle_left_alpha[54][44] = 1'b0; \
	doodle_left_alpha[54][45] = 1'b0; \
	doodle_left_alpha[54][46] = 1'b0; \
	doodle_left_alpha[54][47] = 1'b0; \
	doodle_left_alpha[54][48] = 1'b0; \
	doodle_left_alpha[54][49] = 1'b0; \
	doodle_left_alpha[54][50] = 1'b0; \
	doodle_left_alpha[54][51] = 1'b0; \
	doodle_left_alpha[54][52] = 1'b0; \
	doodle_left_alpha[54][53] = 1'b0; \
	doodle_left_alpha[54][54] = 1'b0; \
	doodle_left_alpha[54][55] = 1'b0; \
	doodle_left_alpha[54][56] = 1'b0; \
	doodle_left_alpha[54][57] = 1'b0; \
	doodle_left_alpha[54][58] = 1'b0; \
	doodle_left_alpha[54][59] = 1'b0; \
	doodle_left_alpha[54][60] = 1'b0; \
	doodle_left_alpha[54][61] = 1'b0; \
	doodle_left_alpha[54][62] = 1'b0; \
	doodle_left_alpha[54][63] = 1'b0; \
	doodle_left_alpha[54][64] = 1'b0; \
	doodle_left_alpha[54][65] = 1'b1; \
	doodle_left_alpha[54][66] = 1'b1; \
	doodle_left_alpha[54][67] = 1'b1; \
	doodle_left_alpha[54][68] = 1'b1; \
	doodle_left_alpha[54][69] = 1'b1; \
	doodle_left_alpha[54][70] = 1'b1; \
	doodle_left_alpha[54][71] = 1'b1; \
	doodle_left_alpha[54][72] = 1'b1; \
	doodle_left_alpha[54][73] = 1'b1; \
	doodle_left_alpha[54][74] = 1'b1; \
	doodle_left_alpha[54][75] = 1'b1; \
	doodle_left_alpha[54][76] = 1'b1; \
	doodle_left_alpha[54][77] = 1'b1; \
	doodle_left_alpha[54][78] = 1'b1; \
	doodle_left_alpha[54][79] = 1'b1; \
	doodle_left_alpha[55][0] = 1'b1; \
	doodle_left_alpha[55][1] = 1'b1; \
	doodle_left_alpha[55][2] = 1'b1; \
	doodle_left_alpha[55][3] = 1'b1; \
	doodle_left_alpha[55][4] = 1'b1; \
	doodle_left_alpha[55][5] = 1'b1; \
	doodle_left_alpha[55][6] = 1'b1; \
	doodle_left_alpha[55][7] = 1'b1; \
	doodle_left_alpha[55][8] = 1'b1; \
	doodle_left_alpha[55][9] = 1'b1; \
	doodle_left_alpha[55][10] = 1'b1; \
	doodle_left_alpha[55][11] = 1'b1; \
	doodle_left_alpha[55][12] = 1'b1; \
	doodle_left_alpha[55][13] = 1'b1; \
	doodle_left_alpha[55][14] = 1'b1; \
	doodle_left_alpha[55][15] = 1'b1; \
	doodle_left_alpha[55][16] = 1'b1; \
	doodle_left_alpha[55][17] = 1'b1; \
	doodle_left_alpha[55][18] = 1'b1; \
	doodle_left_alpha[55][19] = 1'b1; \
	doodle_left_alpha[55][20] = 1'b1; \
	doodle_left_alpha[55][21] = 1'b1; \
	doodle_left_alpha[55][22] = 1'b1; \
	doodle_left_alpha[55][23] = 1'b0; \
	doodle_left_alpha[55][24] = 1'b0; \
	doodle_left_alpha[55][25] = 1'b0; \
	doodle_left_alpha[55][26] = 1'b0; \
	doodle_left_alpha[55][27] = 1'b0; \
	doodle_left_alpha[55][28] = 1'b0; \
	doodle_left_alpha[55][29] = 1'b0; \
	doodle_left_alpha[55][30] = 1'b0; \
	doodle_left_alpha[55][31] = 1'b0; \
	doodle_left_alpha[55][32] = 1'b0; \
	doodle_left_alpha[55][33] = 1'b0; \
	doodle_left_alpha[55][34] = 1'b0; \
	doodle_left_alpha[55][35] = 1'b0; \
	doodle_left_alpha[55][36] = 1'b0; \
	doodle_left_alpha[55][37] = 1'b0; \
	doodle_left_alpha[55][38] = 1'b0; \
	doodle_left_alpha[55][39] = 1'b0; \
	doodle_left_alpha[55][40] = 1'b0; \
	doodle_left_alpha[55][41] = 1'b0; \
	doodle_left_alpha[55][42] = 1'b0; \
	doodle_left_alpha[55][43] = 1'b0; \
	doodle_left_alpha[55][44] = 1'b0; \
	doodle_left_alpha[55][45] = 1'b0; \
	doodle_left_alpha[55][46] = 1'b0; \
	doodle_left_alpha[55][47] = 1'b0; \
	doodle_left_alpha[55][48] = 1'b0; \
	doodle_left_alpha[55][49] = 1'b0; \
	doodle_left_alpha[55][50] = 1'b0; \
	doodle_left_alpha[55][51] = 1'b0; \
	doodle_left_alpha[55][52] = 1'b0; \
	doodle_left_alpha[55][53] = 1'b0; \
	doodle_left_alpha[55][54] = 1'b0; \
	doodle_left_alpha[55][55] = 1'b0; \
	doodle_left_alpha[55][56] = 1'b0; \
	doodle_left_alpha[55][57] = 1'b0; \
	doodle_left_alpha[55][58] = 1'b0; \
	doodle_left_alpha[55][59] = 1'b0; \
	doodle_left_alpha[55][60] = 1'b0; \
	doodle_left_alpha[55][61] = 1'b0; \
	doodle_left_alpha[55][62] = 1'b0; \
	doodle_left_alpha[55][63] = 1'b0; \
	doodle_left_alpha[55][64] = 1'b0; \
	doodle_left_alpha[55][65] = 1'b1; \
	doodle_left_alpha[55][66] = 1'b1; \
	doodle_left_alpha[55][67] = 1'b1; \
	doodle_left_alpha[55][68] = 1'b1; \
	doodle_left_alpha[55][69] = 1'b1; \
	doodle_left_alpha[55][70] = 1'b1; \
	doodle_left_alpha[55][71] = 1'b1; \
	doodle_left_alpha[55][72] = 1'b1; \
	doodle_left_alpha[55][73] = 1'b1; \
	doodle_left_alpha[55][74] = 1'b1; \
	doodle_left_alpha[55][75] = 1'b1; \
	doodle_left_alpha[55][76] = 1'b1; \
	doodle_left_alpha[55][77] = 1'b1; \
	doodle_left_alpha[55][78] = 1'b1; \
	doodle_left_alpha[55][79] = 1'b1; \
	doodle_left_alpha[56][0] = 1'b1; \
	doodle_left_alpha[56][1] = 1'b1; \
	doodle_left_alpha[56][2] = 1'b1; \
	doodle_left_alpha[56][3] = 1'b1; \
	doodle_left_alpha[56][4] = 1'b1; \
	doodle_left_alpha[56][5] = 1'b1; \
	doodle_left_alpha[56][6] = 1'b1; \
	doodle_left_alpha[56][7] = 1'b1; \
	doodle_left_alpha[56][8] = 1'b1; \
	doodle_left_alpha[56][9] = 1'b1; \
	doodle_left_alpha[56][10] = 1'b1; \
	doodle_left_alpha[56][11] = 1'b1; \
	doodle_left_alpha[56][12] = 1'b1; \
	doodle_left_alpha[56][13] = 1'b1; \
	doodle_left_alpha[56][14] = 1'b1; \
	doodle_left_alpha[56][15] = 1'b1; \
	doodle_left_alpha[56][16] = 1'b1; \
	doodle_left_alpha[56][17] = 1'b1; \
	doodle_left_alpha[56][18] = 1'b1; \
	doodle_left_alpha[56][19] = 1'b1; \
	doodle_left_alpha[56][20] = 1'b1; \
	doodle_left_alpha[56][21] = 1'b1; \
	doodle_left_alpha[56][22] = 1'b1; \
	doodle_left_alpha[56][23] = 1'b0; \
	doodle_left_alpha[56][24] = 1'b0; \
	doodle_left_alpha[56][25] = 1'b0; \
	doodle_left_alpha[56][26] = 1'b0; \
	doodle_left_alpha[56][27] = 1'b0; \
	doodle_left_alpha[56][28] = 1'b0; \
	doodle_left_alpha[56][29] = 1'b0; \
	doodle_left_alpha[56][30] = 1'b0; \
	doodle_left_alpha[56][31] = 1'b0; \
	doodle_left_alpha[56][32] = 1'b0; \
	doodle_left_alpha[56][33] = 1'b0; \
	doodle_left_alpha[56][34] = 1'b0; \
	doodle_left_alpha[56][35] = 1'b0; \
	doodle_left_alpha[56][36] = 1'b0; \
	doodle_left_alpha[56][37] = 1'b0; \
	doodle_left_alpha[56][38] = 1'b0; \
	doodle_left_alpha[56][39] = 1'b0; \
	doodle_left_alpha[56][40] = 1'b0; \
	doodle_left_alpha[56][41] = 1'b0; \
	doodle_left_alpha[56][42] = 1'b0; \
	doodle_left_alpha[56][43] = 1'b0; \
	doodle_left_alpha[56][44] = 1'b0; \
	doodle_left_alpha[56][45] = 1'b0; \
	doodle_left_alpha[56][46] = 1'b0; \
	doodle_left_alpha[56][47] = 1'b0; \
	doodle_left_alpha[56][48] = 1'b0; \
	doodle_left_alpha[56][49] = 1'b0; \
	doodle_left_alpha[56][50] = 1'b0; \
	doodle_left_alpha[56][51] = 1'b0; \
	doodle_left_alpha[56][52] = 1'b0; \
	doodle_left_alpha[56][53] = 1'b0; \
	doodle_left_alpha[56][54] = 1'b0; \
	doodle_left_alpha[56][55] = 1'b0; \
	doodle_left_alpha[56][56] = 1'b0; \
	doodle_left_alpha[56][57] = 1'b0; \
	doodle_left_alpha[56][58] = 1'b0; \
	doodle_left_alpha[56][59] = 1'b0; \
	doodle_left_alpha[56][60] = 1'b0; \
	doodle_left_alpha[56][61] = 1'b0; \
	doodle_left_alpha[56][62] = 1'b0; \
	doodle_left_alpha[56][63] = 1'b0; \
	doodle_left_alpha[56][64] = 1'b0; \
	doodle_left_alpha[56][65] = 1'b1; \
	doodle_left_alpha[56][66] = 1'b1; \
	doodle_left_alpha[56][67] = 1'b1; \
	doodle_left_alpha[56][68] = 1'b1; \
	doodle_left_alpha[56][69] = 1'b1; \
	doodle_left_alpha[56][70] = 1'b1; \
	doodle_left_alpha[56][71] = 1'b1; \
	doodle_left_alpha[56][72] = 1'b1; \
	doodle_left_alpha[56][73] = 1'b1; \
	doodle_left_alpha[56][74] = 1'b1; \
	doodle_left_alpha[56][75] = 1'b1; \
	doodle_left_alpha[56][76] = 1'b1; \
	doodle_left_alpha[56][77] = 1'b1; \
	doodle_left_alpha[56][78] = 1'b1; \
	doodle_left_alpha[56][79] = 1'b1; \
	doodle_left_alpha[57][0] = 1'b1; \
	doodle_left_alpha[57][1] = 1'b1; \
	doodle_left_alpha[57][2] = 1'b1; \
	doodle_left_alpha[57][3] = 1'b1; \
	doodle_left_alpha[57][4] = 1'b1; \
	doodle_left_alpha[57][5] = 1'b1; \
	doodle_left_alpha[57][6] = 1'b1; \
	doodle_left_alpha[57][7] = 1'b1; \
	doodle_left_alpha[57][8] = 1'b1; \
	doodle_left_alpha[57][9] = 1'b1; \
	doodle_left_alpha[57][10] = 1'b1; \
	doodle_left_alpha[57][11] = 1'b1; \
	doodle_left_alpha[57][12] = 1'b1; \
	doodle_left_alpha[57][13] = 1'b1; \
	doodle_left_alpha[57][14] = 1'b1; \
	doodle_left_alpha[57][15] = 1'b1; \
	doodle_left_alpha[57][16] = 1'b1; \
	doodle_left_alpha[57][17] = 1'b1; \
	doodle_left_alpha[57][18] = 1'b1; \
	doodle_left_alpha[57][19] = 1'b1; \
	doodle_left_alpha[57][20] = 1'b1; \
	doodle_left_alpha[57][21] = 1'b1; \
	doodle_left_alpha[57][22] = 1'b1; \
	doodle_left_alpha[57][23] = 1'b0; \
	doodle_left_alpha[57][24] = 1'b0; \
	doodle_left_alpha[57][25] = 1'b0; \
	doodle_left_alpha[57][26] = 1'b0; \
	doodle_left_alpha[57][27] = 1'b0; \
	doodle_left_alpha[57][28] = 1'b0; \
	doodle_left_alpha[57][29] = 1'b0; \
	doodle_left_alpha[57][30] = 1'b0; \
	doodle_left_alpha[57][31] = 1'b0; \
	doodle_left_alpha[57][32] = 1'b0; \
	doodle_left_alpha[57][33] = 1'b0; \
	doodle_left_alpha[57][34] = 1'b0; \
	doodle_left_alpha[57][35] = 1'b0; \
	doodle_left_alpha[57][36] = 1'b0; \
	doodle_left_alpha[57][37] = 1'b0; \
	doodle_left_alpha[57][38] = 1'b0; \
	doodle_left_alpha[57][39] = 1'b0; \
	doodle_left_alpha[57][40] = 1'b0; \
	doodle_left_alpha[57][41] = 1'b0; \
	doodle_left_alpha[57][42] = 1'b0; \
	doodle_left_alpha[57][43] = 1'b0; \
	doodle_left_alpha[57][44] = 1'b0; \
	doodle_left_alpha[57][45] = 1'b0; \
	doodle_left_alpha[57][46] = 1'b0; \
	doodle_left_alpha[57][47] = 1'b0; \
	doodle_left_alpha[57][48] = 1'b0; \
	doodle_left_alpha[57][49] = 1'b0; \
	doodle_left_alpha[57][50] = 1'b0; \
	doodle_left_alpha[57][51] = 1'b0; \
	doodle_left_alpha[57][52] = 1'b0; \
	doodle_left_alpha[57][53] = 1'b0; \
	doodle_left_alpha[57][54] = 1'b0; \
	doodle_left_alpha[57][55] = 1'b0; \
	doodle_left_alpha[57][56] = 1'b0; \
	doodle_left_alpha[57][57] = 1'b0; \
	doodle_left_alpha[57][58] = 1'b0; \
	doodle_left_alpha[57][59] = 1'b0; \
	doodle_left_alpha[57][60] = 1'b0; \
	doodle_left_alpha[57][61] = 1'b0; \
	doodle_left_alpha[57][62] = 1'b0; \
	doodle_left_alpha[57][63] = 1'b0; \
	doodle_left_alpha[57][64] = 1'b0; \
	doodle_left_alpha[57][65] = 1'b1; \
	doodle_left_alpha[57][66] = 1'b1; \
	doodle_left_alpha[57][67] = 1'b1; \
	doodle_left_alpha[57][68] = 1'b1; \
	doodle_left_alpha[57][69] = 1'b1; \
	doodle_left_alpha[57][70] = 1'b1; \
	doodle_left_alpha[57][71] = 1'b1; \
	doodle_left_alpha[57][72] = 1'b1; \
	doodle_left_alpha[57][73] = 1'b1; \
	doodle_left_alpha[57][74] = 1'b1; \
	doodle_left_alpha[57][75] = 1'b1; \
	doodle_left_alpha[57][76] = 1'b1; \
	doodle_left_alpha[57][77] = 1'b1; \
	doodle_left_alpha[57][78] = 1'b1; \
	doodle_left_alpha[57][79] = 1'b1; \
	doodle_left_alpha[58][0] = 1'b1; \
	doodle_left_alpha[58][1] = 1'b1; \
	doodle_left_alpha[58][2] = 1'b1; \
	doodle_left_alpha[58][3] = 1'b1; \
	doodle_left_alpha[58][4] = 1'b1; \
	doodle_left_alpha[58][5] = 1'b1; \
	doodle_left_alpha[58][6] = 1'b1; \
	doodle_left_alpha[58][7] = 1'b1; \
	doodle_left_alpha[58][8] = 1'b1; \
	doodle_left_alpha[58][9] = 1'b1; \
	doodle_left_alpha[58][10] = 1'b1; \
	doodle_left_alpha[58][11] = 1'b1; \
	doodle_left_alpha[58][12] = 1'b1; \
	doodle_left_alpha[58][13] = 1'b1; \
	doodle_left_alpha[58][14] = 1'b1; \
	doodle_left_alpha[58][15] = 1'b1; \
	doodle_left_alpha[58][16] = 1'b1; \
	doodle_left_alpha[58][17] = 1'b1; \
	doodle_left_alpha[58][18] = 1'b1; \
	doodle_left_alpha[58][19] = 1'b1; \
	doodle_left_alpha[58][20] = 1'b1; \
	doodle_left_alpha[58][21] = 1'b1; \
	doodle_left_alpha[58][22] = 1'b1; \
	doodle_left_alpha[58][23] = 1'b0; \
	doodle_left_alpha[58][24] = 1'b0; \
	doodle_left_alpha[58][25] = 1'b0; \
	doodle_left_alpha[58][26] = 1'b0; \
	doodle_left_alpha[58][27] = 1'b0; \
	doodle_left_alpha[58][28] = 1'b0; \
	doodle_left_alpha[58][29] = 1'b0; \
	doodle_left_alpha[58][30] = 1'b0; \
	doodle_left_alpha[58][31] = 1'b0; \
	doodle_left_alpha[58][32] = 1'b0; \
	doodle_left_alpha[58][33] = 1'b0; \
	doodle_left_alpha[58][34] = 1'b0; \
	doodle_left_alpha[58][35] = 1'b0; \
	doodle_left_alpha[58][36] = 1'b0; \
	doodle_left_alpha[58][37] = 1'b0; \
	doodle_left_alpha[58][38] = 1'b0; \
	doodle_left_alpha[58][39] = 1'b0; \
	doodle_left_alpha[58][40] = 1'b0; \
	doodle_left_alpha[58][41] = 1'b0; \
	doodle_left_alpha[58][42] = 1'b0; \
	doodle_left_alpha[58][43] = 1'b0; \
	doodle_left_alpha[58][44] = 1'b0; \
	doodle_left_alpha[58][45] = 1'b0; \
	doodle_left_alpha[58][46] = 1'b0; \
	doodle_left_alpha[58][47] = 1'b0; \
	doodle_left_alpha[58][48] = 1'b0; \
	doodle_left_alpha[58][49] = 1'b0; \
	doodle_left_alpha[58][50] = 1'b0; \
	doodle_left_alpha[58][51] = 1'b0; \
	doodle_left_alpha[58][52] = 1'b0; \
	doodle_left_alpha[58][53] = 1'b0; \
	doodle_left_alpha[58][54] = 1'b0; \
	doodle_left_alpha[58][55] = 1'b0; \
	doodle_left_alpha[58][56] = 1'b0; \
	doodle_left_alpha[58][57] = 1'b0; \
	doodle_left_alpha[58][58] = 1'b0; \
	doodle_left_alpha[58][59] = 1'b0; \
	doodle_left_alpha[58][60] = 1'b0; \
	doodle_left_alpha[58][61] = 1'b0; \
	doodle_left_alpha[58][62] = 1'b0; \
	doodle_left_alpha[58][63] = 1'b0; \
	doodle_left_alpha[58][64] = 1'b0; \
	doodle_left_alpha[58][65] = 1'b1; \
	doodle_left_alpha[58][66] = 1'b1; \
	doodle_left_alpha[58][67] = 1'b1; \
	doodle_left_alpha[58][68] = 1'b1; \
	doodle_left_alpha[58][69] = 1'b1; \
	doodle_left_alpha[58][70] = 1'b1; \
	doodle_left_alpha[58][71] = 1'b1; \
	doodle_left_alpha[58][72] = 1'b1; \
	doodle_left_alpha[58][73] = 1'b1; \
	doodle_left_alpha[58][74] = 1'b1; \
	doodle_left_alpha[58][75] = 1'b1; \
	doodle_left_alpha[58][76] = 1'b1; \
	doodle_left_alpha[58][77] = 1'b1; \
	doodle_left_alpha[58][78] = 1'b1; \
	doodle_left_alpha[58][79] = 1'b1; \
	doodle_left_alpha[59][0] = 1'b1; \
	doodle_left_alpha[59][1] = 1'b1; \
	doodle_left_alpha[59][2] = 1'b1; \
	doodle_left_alpha[59][3] = 1'b1; \
	doodle_left_alpha[59][4] = 1'b1; \
	doodle_left_alpha[59][5] = 1'b1; \
	doodle_left_alpha[59][6] = 1'b1; \
	doodle_left_alpha[59][7] = 1'b1; \
	doodle_left_alpha[59][8] = 1'b1; \
	doodle_left_alpha[59][9] = 1'b1; \
	doodle_left_alpha[59][10] = 1'b1; \
	doodle_left_alpha[59][11] = 1'b1; \
	doodle_left_alpha[59][12] = 1'b1; \
	doodle_left_alpha[59][13] = 1'b1; \
	doodle_left_alpha[59][14] = 1'b1; \
	doodle_left_alpha[59][15] = 1'b1; \
	doodle_left_alpha[59][16] = 1'b1; \
	doodle_left_alpha[59][17] = 1'b1; \
	doodle_left_alpha[59][18] = 1'b1; \
	doodle_left_alpha[59][19] = 1'b1; \
	doodle_left_alpha[59][20] = 1'b1; \
	doodle_left_alpha[59][21] = 1'b1; \
	doodle_left_alpha[59][22] = 1'b1; \
	doodle_left_alpha[59][23] = 1'b0; \
	doodle_left_alpha[59][24] = 1'b0; \
	doodle_left_alpha[59][25] = 1'b0; \
	doodle_left_alpha[59][26] = 1'b0; \
	doodle_left_alpha[59][27] = 1'b0; \
	doodle_left_alpha[59][28] = 1'b0; \
	doodle_left_alpha[59][29] = 1'b0; \
	doodle_left_alpha[59][30] = 1'b0; \
	doodle_left_alpha[59][31] = 1'b0; \
	doodle_left_alpha[59][32] = 1'b0; \
	doodle_left_alpha[59][33] = 1'b0; \
	doodle_left_alpha[59][34] = 1'b0; \
	doodle_left_alpha[59][35] = 1'b0; \
	doodle_left_alpha[59][36] = 1'b0; \
	doodle_left_alpha[59][37] = 1'b0; \
	doodle_left_alpha[59][38] = 1'b0; \
	doodle_left_alpha[59][39] = 1'b0; \
	doodle_left_alpha[59][40] = 1'b0; \
	doodle_left_alpha[59][41] = 1'b0; \
	doodle_left_alpha[59][42] = 1'b0; \
	doodle_left_alpha[59][43] = 1'b0; \
	doodle_left_alpha[59][44] = 1'b0; \
	doodle_left_alpha[59][45] = 1'b0; \
	doodle_left_alpha[59][46] = 1'b0; \
	doodle_left_alpha[59][47] = 1'b0; \
	doodle_left_alpha[59][48] = 1'b0; \
	doodle_left_alpha[59][49] = 1'b0; \
	doodle_left_alpha[59][50] = 1'b0; \
	doodle_left_alpha[59][51] = 1'b0; \
	doodle_left_alpha[59][52] = 1'b0; \
	doodle_left_alpha[59][53] = 1'b0; \
	doodle_left_alpha[59][54] = 1'b0; \
	doodle_left_alpha[59][55] = 1'b0; \
	doodle_left_alpha[59][56] = 1'b0; \
	doodle_left_alpha[59][57] = 1'b0; \
	doodle_left_alpha[59][58] = 1'b0; \
	doodle_left_alpha[59][59] = 1'b0; \
	doodle_left_alpha[59][60] = 1'b0; \
	doodle_left_alpha[59][61] = 1'b0; \
	doodle_left_alpha[59][62] = 1'b0; \
	doodle_left_alpha[59][63] = 1'b0; \
	doodle_left_alpha[59][64] = 1'b0; \
	doodle_left_alpha[59][65] = 1'b1; \
	doodle_left_alpha[59][66] = 1'b1; \
	doodle_left_alpha[59][67] = 1'b1; \
	doodle_left_alpha[59][68] = 1'b1; \
	doodle_left_alpha[59][69] = 1'b1; \
	doodle_left_alpha[59][70] = 1'b1; \
	doodle_left_alpha[59][71] = 1'b1; \
	doodle_left_alpha[59][72] = 1'b1; \
	doodle_left_alpha[59][73] = 1'b1; \
	doodle_left_alpha[59][74] = 1'b1; \
	doodle_left_alpha[59][75] = 1'b1; \
	doodle_left_alpha[59][76] = 1'b1; \
	doodle_left_alpha[59][77] = 1'b1; \
	doodle_left_alpha[59][78] = 1'b1; \
	doodle_left_alpha[59][79] = 1'b1; \
	doodle_left_alpha[60][0] = 1'b1; \
	doodle_left_alpha[60][1] = 1'b1; \
	doodle_left_alpha[60][2] = 1'b1; \
	doodle_left_alpha[60][3] = 1'b1; \
	doodle_left_alpha[60][4] = 1'b1; \
	doodle_left_alpha[60][5] = 1'b1; \
	doodle_left_alpha[60][6] = 1'b1; \
	doodle_left_alpha[60][7] = 1'b1; \
	doodle_left_alpha[60][8] = 1'b1; \
	doodle_left_alpha[60][9] = 1'b1; \
	doodle_left_alpha[60][10] = 1'b1; \
	doodle_left_alpha[60][11] = 1'b1; \
	doodle_left_alpha[60][12] = 1'b1; \
	doodle_left_alpha[60][13] = 1'b1; \
	doodle_left_alpha[60][14] = 1'b1; \
	doodle_left_alpha[60][15] = 1'b1; \
	doodle_left_alpha[60][16] = 1'b1; \
	doodle_left_alpha[60][17] = 1'b1; \
	doodle_left_alpha[60][18] = 1'b1; \
	doodle_left_alpha[60][19] = 1'b1; \
	doodle_left_alpha[60][20] = 1'b1; \
	doodle_left_alpha[60][21] = 1'b1; \
	doodle_left_alpha[60][22] = 1'b1; \
	doodle_left_alpha[60][23] = 1'b0; \
	doodle_left_alpha[60][24] = 1'b0; \
	doodle_left_alpha[60][25] = 1'b0; \
	doodle_left_alpha[60][26] = 1'b0; \
	doodle_left_alpha[60][27] = 1'b0; \
	doodle_left_alpha[60][28] = 1'b0; \
	doodle_left_alpha[60][29] = 1'b0; \
	doodle_left_alpha[60][30] = 1'b0; \
	doodle_left_alpha[60][31] = 1'b0; \
	doodle_left_alpha[60][32] = 1'b0; \
	doodle_left_alpha[60][33] = 1'b0; \
	doodle_left_alpha[60][34] = 1'b0; \
	doodle_left_alpha[60][35] = 1'b0; \
	doodle_left_alpha[60][36] = 1'b0; \
	doodle_left_alpha[60][37] = 1'b0; \
	doodle_left_alpha[60][38] = 1'b0; \
	doodle_left_alpha[60][39] = 1'b0; \
	doodle_left_alpha[60][40] = 1'b0; \
	doodle_left_alpha[60][41] = 1'b0; \
	doodle_left_alpha[60][42] = 1'b0; \
	doodle_left_alpha[60][43] = 1'b0; \
	doodle_left_alpha[60][44] = 1'b0; \
	doodle_left_alpha[60][45] = 1'b0; \
	doodle_left_alpha[60][46] = 1'b0; \
	doodle_left_alpha[60][47] = 1'b0; \
	doodle_left_alpha[60][48] = 1'b0; \
	doodle_left_alpha[60][49] = 1'b0; \
	doodle_left_alpha[60][50] = 1'b0; \
	doodle_left_alpha[60][51] = 1'b0; \
	doodle_left_alpha[60][52] = 1'b0; \
	doodle_left_alpha[60][53] = 1'b0; \
	doodle_left_alpha[60][54] = 1'b0; \
	doodle_left_alpha[60][55] = 1'b0; \
	doodle_left_alpha[60][56] = 1'b0; \
	doodle_left_alpha[60][57] = 1'b0; \
	doodle_left_alpha[60][58] = 1'b0; \
	doodle_left_alpha[60][59] = 1'b0; \
	doodle_left_alpha[60][60] = 1'b0; \
	doodle_left_alpha[60][61] = 1'b0; \
	doodle_left_alpha[60][62] = 1'b0; \
	doodle_left_alpha[60][63] = 1'b0; \
	doodle_left_alpha[60][64] = 1'b0; \
	doodle_left_alpha[60][65] = 1'b1; \
	doodle_left_alpha[60][66] = 1'b1; \
	doodle_left_alpha[60][67] = 1'b1; \
	doodle_left_alpha[60][68] = 1'b1; \
	doodle_left_alpha[60][69] = 1'b1; \
	doodle_left_alpha[60][70] = 1'b1; \
	doodle_left_alpha[60][71] = 1'b1; \
	doodle_left_alpha[60][72] = 1'b1; \
	doodle_left_alpha[60][73] = 1'b1; \
	doodle_left_alpha[60][74] = 1'b1; \
	doodle_left_alpha[60][75] = 1'b1; \
	doodle_left_alpha[60][76] = 1'b1; \
	doodle_left_alpha[60][77] = 1'b1; \
	doodle_left_alpha[60][78] = 1'b1; \
	doodle_left_alpha[60][79] = 1'b1; \
	doodle_left_alpha[61][0] = 1'b1; \
	doodle_left_alpha[61][1] = 1'b1; \
	doodle_left_alpha[61][2] = 1'b1; \
	doodle_left_alpha[61][3] = 1'b1; \
	doodle_left_alpha[61][4] = 1'b1; \
	doodle_left_alpha[61][5] = 1'b1; \
	doodle_left_alpha[61][6] = 1'b1; \
	doodle_left_alpha[61][7] = 1'b1; \
	doodle_left_alpha[61][8] = 1'b1; \
	doodle_left_alpha[61][9] = 1'b1; \
	doodle_left_alpha[61][10] = 1'b1; \
	doodle_left_alpha[61][11] = 1'b1; \
	doodle_left_alpha[61][12] = 1'b1; \
	doodle_left_alpha[61][13] = 1'b1; \
	doodle_left_alpha[61][14] = 1'b1; \
	doodle_left_alpha[61][15] = 1'b1; \
	doodle_left_alpha[61][16] = 1'b1; \
	doodle_left_alpha[61][17] = 1'b1; \
	doodle_left_alpha[61][18] = 1'b1; \
	doodle_left_alpha[61][19] = 1'b1; \
	doodle_left_alpha[61][20] = 1'b1; \
	doodle_left_alpha[61][21] = 1'b1; \
	doodle_left_alpha[61][22] = 1'b1; \
	doodle_left_alpha[61][23] = 1'b0; \
	doodle_left_alpha[61][24] = 1'b0; \
	doodle_left_alpha[61][25] = 1'b0; \
	doodle_left_alpha[61][26] = 1'b0; \
	doodle_left_alpha[61][27] = 1'b0; \
	doodle_left_alpha[61][28] = 1'b0; \
	doodle_left_alpha[61][29] = 1'b0; \
	doodle_left_alpha[61][30] = 1'b0; \
	doodle_left_alpha[61][31] = 1'b0; \
	doodle_left_alpha[61][32] = 1'b0; \
	doodle_left_alpha[61][33] = 1'b0; \
	doodle_left_alpha[61][34] = 1'b0; \
	doodle_left_alpha[61][35] = 1'b0; \
	doodle_left_alpha[61][36] = 1'b0; \
	doodle_left_alpha[61][37] = 1'b0; \
	doodle_left_alpha[61][38] = 1'b0; \
	doodle_left_alpha[61][39] = 1'b0; \
	doodle_left_alpha[61][40] = 1'b0; \
	doodle_left_alpha[61][41] = 1'b0; \
	doodle_left_alpha[61][42] = 1'b0; \
	doodle_left_alpha[61][43] = 1'b0; \
	doodle_left_alpha[61][44] = 1'b0; \
	doodle_left_alpha[61][45] = 1'b0; \
	doodle_left_alpha[61][46] = 1'b0; \
	doodle_left_alpha[61][47] = 1'b0; \
	doodle_left_alpha[61][48] = 1'b0; \
	doodle_left_alpha[61][49] = 1'b0; \
	doodle_left_alpha[61][50] = 1'b0; \
	doodle_left_alpha[61][51] = 1'b0; \
	doodle_left_alpha[61][52] = 1'b0; \
	doodle_left_alpha[61][53] = 1'b0; \
	doodle_left_alpha[61][54] = 1'b0; \
	doodle_left_alpha[61][55] = 1'b0; \
	doodle_left_alpha[61][56] = 1'b0; \
	doodle_left_alpha[61][57] = 1'b0; \
	doodle_left_alpha[61][58] = 1'b0; \
	doodle_left_alpha[61][59] = 1'b0; \
	doodle_left_alpha[61][60] = 1'b0; \
	doodle_left_alpha[61][61] = 1'b0; \
	doodle_left_alpha[61][62] = 1'b0; \
	doodle_left_alpha[61][63] = 1'b0; \
	doodle_left_alpha[61][64] = 1'b0; \
	doodle_left_alpha[61][65] = 1'b1; \
	doodle_left_alpha[61][66] = 1'b1; \
	doodle_left_alpha[61][67] = 1'b1; \
	doodle_left_alpha[61][68] = 1'b1; \
	doodle_left_alpha[61][69] = 1'b1; \
	doodle_left_alpha[61][70] = 1'b1; \
	doodle_left_alpha[61][71] = 1'b1; \
	doodle_left_alpha[61][72] = 1'b1; \
	doodle_left_alpha[61][73] = 1'b1; \
	doodle_left_alpha[61][74] = 1'b1; \
	doodle_left_alpha[61][75] = 1'b1; \
	doodle_left_alpha[61][76] = 1'b1; \
	doodle_left_alpha[61][77] = 1'b1; \
	doodle_left_alpha[61][78] = 1'b1; \
	doodle_left_alpha[61][79] = 1'b1; \
	doodle_left_alpha[62][0] = 1'b1; \
	doodle_left_alpha[62][1] = 1'b1; \
	doodle_left_alpha[62][2] = 1'b1; \
	doodle_left_alpha[62][3] = 1'b1; \
	doodle_left_alpha[62][4] = 1'b1; \
	doodle_left_alpha[62][5] = 1'b1; \
	doodle_left_alpha[62][6] = 1'b1; \
	doodle_left_alpha[62][7] = 1'b1; \
	doodle_left_alpha[62][8] = 1'b1; \
	doodle_left_alpha[62][9] = 1'b1; \
	doodle_left_alpha[62][10] = 1'b1; \
	doodle_left_alpha[62][11] = 1'b1; \
	doodle_left_alpha[62][12] = 1'b1; \
	doodle_left_alpha[62][13] = 1'b1; \
	doodle_left_alpha[62][14] = 1'b1; \
	doodle_left_alpha[62][15] = 1'b1; \
	doodle_left_alpha[62][16] = 1'b1; \
	doodle_left_alpha[62][17] = 1'b1; \
	doodle_left_alpha[62][18] = 1'b1; \
	doodle_left_alpha[62][19] = 1'b1; \
	doodle_left_alpha[62][20] = 1'b1; \
	doodle_left_alpha[62][21] = 1'b1; \
	doodle_left_alpha[62][22] = 1'b1; \
	doodle_left_alpha[62][23] = 1'b0; \
	doodle_left_alpha[62][24] = 1'b0; \
	doodle_left_alpha[62][25] = 1'b0; \
	doodle_left_alpha[62][26] = 1'b0; \
	doodle_left_alpha[62][27] = 1'b0; \
	doodle_left_alpha[62][28] = 1'b0; \
	doodle_left_alpha[62][29] = 1'b0; \
	doodle_left_alpha[62][30] = 1'b0; \
	doodle_left_alpha[62][31] = 1'b0; \
	doodle_left_alpha[62][32] = 1'b0; \
	doodle_left_alpha[62][33] = 1'b0; \
	doodle_left_alpha[62][34] = 1'b0; \
	doodle_left_alpha[62][35] = 1'b0; \
	doodle_left_alpha[62][36] = 1'b0; \
	doodle_left_alpha[62][37] = 1'b0; \
	doodle_left_alpha[62][38] = 1'b0; \
	doodle_left_alpha[62][39] = 1'b0; \
	doodle_left_alpha[62][40] = 1'b0; \
	doodle_left_alpha[62][41] = 1'b0; \
	doodle_left_alpha[62][42] = 1'b0; \
	doodle_left_alpha[62][43] = 1'b0; \
	doodle_left_alpha[62][44] = 1'b0; \
	doodle_left_alpha[62][45] = 1'b0; \
	doodle_left_alpha[62][46] = 1'b0; \
	doodle_left_alpha[62][47] = 1'b0; \
	doodle_left_alpha[62][48] = 1'b0; \
	doodle_left_alpha[62][49] = 1'b0; \
	doodle_left_alpha[62][50] = 1'b0; \
	doodle_left_alpha[62][51] = 1'b0; \
	doodle_left_alpha[62][52] = 1'b0; \
	doodle_left_alpha[62][53] = 1'b0; \
	doodle_left_alpha[62][54] = 1'b0; \
	doodle_left_alpha[62][55] = 1'b0; \
	doodle_left_alpha[62][56] = 1'b0; \
	doodle_left_alpha[62][57] = 1'b0; \
	doodle_left_alpha[62][58] = 1'b0; \
	doodle_left_alpha[62][59] = 1'b0; \
	doodle_left_alpha[62][60] = 1'b0; \
	doodle_left_alpha[62][61] = 1'b0; \
	doodle_left_alpha[62][62] = 1'b0; \
	doodle_left_alpha[62][63] = 1'b0; \
	doodle_left_alpha[62][64] = 1'b0; \
	doodle_left_alpha[62][65] = 1'b1; \
	doodle_left_alpha[62][66] = 1'b1; \
	doodle_left_alpha[62][67] = 1'b1; \
	doodle_left_alpha[62][68] = 1'b1; \
	doodle_left_alpha[62][69] = 1'b1; \
	doodle_left_alpha[62][70] = 1'b1; \
	doodle_left_alpha[62][71] = 1'b1; \
	doodle_left_alpha[62][72] = 1'b1; \
	doodle_left_alpha[62][73] = 1'b1; \
	doodle_left_alpha[62][74] = 1'b1; \
	doodle_left_alpha[62][75] = 1'b1; \
	doodle_left_alpha[62][76] = 1'b1; \
	doodle_left_alpha[62][77] = 1'b1; \
	doodle_left_alpha[62][78] = 1'b1; \
	doodle_left_alpha[62][79] = 1'b1; \
	doodle_left_alpha[63][0] = 1'b1; \
	doodle_left_alpha[63][1] = 1'b1; \
	doodle_left_alpha[63][2] = 1'b1; \
	doodle_left_alpha[63][3] = 1'b1; \
	doodle_left_alpha[63][4] = 1'b1; \
	doodle_left_alpha[63][5] = 1'b1; \
	doodle_left_alpha[63][6] = 1'b1; \
	doodle_left_alpha[63][7] = 1'b1; \
	doodle_left_alpha[63][8] = 1'b1; \
	doodle_left_alpha[63][9] = 1'b1; \
	doodle_left_alpha[63][10] = 1'b1; \
	doodle_left_alpha[63][11] = 1'b1; \
	doodle_left_alpha[63][12] = 1'b1; \
	doodle_left_alpha[63][13] = 1'b1; \
	doodle_left_alpha[63][14] = 1'b1; \
	doodle_left_alpha[63][15] = 1'b1; \
	doodle_left_alpha[63][16] = 1'b1; \
	doodle_left_alpha[63][17] = 1'b1; \
	doodle_left_alpha[63][18] = 1'b1; \
	doodle_left_alpha[63][19] = 1'b1; \
	doodle_left_alpha[63][20] = 1'b1; \
	doodle_left_alpha[63][21] = 1'b1; \
	doodle_left_alpha[63][22] = 1'b1; \
	doodle_left_alpha[63][23] = 1'b0; \
	doodle_left_alpha[63][24] = 1'b0; \
	doodle_left_alpha[63][25] = 1'b0; \
	doodle_left_alpha[63][26] = 1'b0; \
	doodle_left_alpha[63][27] = 1'b0; \
	doodle_left_alpha[63][28] = 1'b0; \
	doodle_left_alpha[63][29] = 1'b0; \
	doodle_left_alpha[63][30] = 1'b0; \
	doodle_left_alpha[63][31] = 1'b0; \
	doodle_left_alpha[63][32] = 1'b0; \
	doodle_left_alpha[63][33] = 1'b0; \
	doodle_left_alpha[63][34] = 1'b0; \
	doodle_left_alpha[63][35] = 1'b0; \
	doodle_left_alpha[63][36] = 1'b0; \
	doodle_left_alpha[63][37] = 1'b0; \
	doodle_left_alpha[63][38] = 1'b0; \
	doodle_left_alpha[63][39] = 1'b0; \
	doodle_left_alpha[63][40] = 1'b0; \
	doodle_left_alpha[63][41] = 1'b0; \
	doodle_left_alpha[63][42] = 1'b0; \
	doodle_left_alpha[63][43] = 1'b0; \
	doodle_left_alpha[63][44] = 1'b0; \
	doodle_left_alpha[63][45] = 1'b0; \
	doodle_left_alpha[63][46] = 1'b0; \
	doodle_left_alpha[63][47] = 1'b0; \
	doodle_left_alpha[63][48] = 1'b0; \
	doodle_left_alpha[63][49] = 1'b0; \
	doodle_left_alpha[63][50] = 1'b0; \
	doodle_left_alpha[63][51] = 1'b0; \
	doodle_left_alpha[63][52] = 1'b0; \
	doodle_left_alpha[63][53] = 1'b0; \
	doodle_left_alpha[63][54] = 1'b0; \
	doodle_left_alpha[63][55] = 1'b0; \
	doodle_left_alpha[63][56] = 1'b0; \
	doodle_left_alpha[63][57] = 1'b0; \
	doodle_left_alpha[63][58] = 1'b0; \
	doodle_left_alpha[63][59] = 1'b0; \
	doodle_left_alpha[63][60] = 1'b0; \
	doodle_left_alpha[63][61] = 1'b0; \
	doodle_left_alpha[63][62] = 1'b0; \
	doodle_left_alpha[63][63] = 1'b0; \
	doodle_left_alpha[63][64] = 1'b0; \
	doodle_left_alpha[63][65] = 1'b1; \
	doodle_left_alpha[63][66] = 1'b1; \
	doodle_left_alpha[63][67] = 1'b1; \
	doodle_left_alpha[63][68] = 1'b1; \
	doodle_left_alpha[63][69] = 1'b1; \
	doodle_left_alpha[63][70] = 1'b1; \
	doodle_left_alpha[63][71] = 1'b1; \
	doodle_left_alpha[63][72] = 1'b1; \
	doodle_left_alpha[63][73] = 1'b1; \
	doodle_left_alpha[63][74] = 1'b1; \
	doodle_left_alpha[63][75] = 1'b1; \
	doodle_left_alpha[63][76] = 1'b1; \
	doodle_left_alpha[63][77] = 1'b1; \
	doodle_left_alpha[63][78] = 1'b1; \
	doodle_left_alpha[63][79] = 1'b1; \
	doodle_left_alpha[64][0] = 1'b1; \
	doodle_left_alpha[64][1] = 1'b1; \
	doodle_left_alpha[64][2] = 1'b1; \
	doodle_left_alpha[64][3] = 1'b1; \
	doodle_left_alpha[64][4] = 1'b1; \
	doodle_left_alpha[64][5] = 1'b1; \
	doodle_left_alpha[64][6] = 1'b1; \
	doodle_left_alpha[64][7] = 1'b1; \
	doodle_left_alpha[64][8] = 1'b1; \
	doodle_left_alpha[64][9] = 1'b1; \
	doodle_left_alpha[64][10] = 1'b1; \
	doodle_left_alpha[64][11] = 1'b1; \
	doodle_left_alpha[64][12] = 1'b1; \
	doodle_left_alpha[64][13] = 1'b1; \
	doodle_left_alpha[64][14] = 1'b1; \
	doodle_left_alpha[64][15] = 1'b1; \
	doodle_left_alpha[64][16] = 1'b1; \
	doodle_left_alpha[64][17] = 1'b1; \
	doodle_left_alpha[64][18] = 1'b1; \
	doodle_left_alpha[64][19] = 1'b1; \
	doodle_left_alpha[64][20] = 1'b1; \
	doodle_left_alpha[64][21] = 1'b1; \
	doodle_left_alpha[64][22] = 1'b1; \
	doodle_left_alpha[64][23] = 1'b0; \
	doodle_left_alpha[64][24] = 1'b0; \
	doodle_left_alpha[64][25] = 1'b0; \
	doodle_left_alpha[64][26] = 1'b0; \
	doodle_left_alpha[64][27] = 1'b0; \
	doodle_left_alpha[64][28] = 1'b0; \
	doodle_left_alpha[64][29] = 1'b0; \
	doodle_left_alpha[64][30] = 1'b0; \
	doodle_left_alpha[64][31] = 1'b0; \
	doodle_left_alpha[64][32] = 1'b0; \
	doodle_left_alpha[64][33] = 1'b0; \
	doodle_left_alpha[64][34] = 1'b0; \
	doodle_left_alpha[64][35] = 1'b0; \
	doodle_left_alpha[64][36] = 1'b0; \
	doodle_left_alpha[64][37] = 1'b0; \
	doodle_left_alpha[64][38] = 1'b0; \
	doodle_left_alpha[64][39] = 1'b0; \
	doodle_left_alpha[64][40] = 1'b0; \
	doodle_left_alpha[64][41] = 1'b0; \
	doodle_left_alpha[64][42] = 1'b0; \
	doodle_left_alpha[64][43] = 1'b0; \
	doodle_left_alpha[64][44] = 1'b0; \
	doodle_left_alpha[64][45] = 1'b0; \
	doodle_left_alpha[64][46] = 1'b0; \
	doodle_left_alpha[64][47] = 1'b0; \
	doodle_left_alpha[64][48] = 1'b0; \
	doodle_left_alpha[64][49] = 1'b0; \
	doodle_left_alpha[64][50] = 1'b0; \
	doodle_left_alpha[64][51] = 1'b0; \
	doodle_left_alpha[64][52] = 1'b0; \
	doodle_left_alpha[64][53] = 1'b0; \
	doodle_left_alpha[64][54] = 1'b0; \
	doodle_left_alpha[64][55] = 1'b0; \
	doodle_left_alpha[64][56] = 1'b0; \
	doodle_left_alpha[64][57] = 1'b0; \
	doodle_left_alpha[64][58] = 1'b0; \
	doodle_left_alpha[64][59] = 1'b0; \
	doodle_left_alpha[64][60] = 1'b0; \
	doodle_left_alpha[64][61] = 1'b0; \
	doodle_left_alpha[64][62] = 1'b0; \
	doodle_left_alpha[64][63] = 1'b0; \
	doodle_left_alpha[64][64] = 1'b0; \
	doodle_left_alpha[64][65] = 1'b1; \
	doodle_left_alpha[64][66] = 1'b1; \
	doodle_left_alpha[64][67] = 1'b1; \
	doodle_left_alpha[64][68] = 1'b1; \
	doodle_left_alpha[64][69] = 1'b1; \
	doodle_left_alpha[64][70] = 1'b1; \
	doodle_left_alpha[64][71] = 1'b1; \
	doodle_left_alpha[64][72] = 1'b1; \
	doodle_left_alpha[64][73] = 1'b1; \
	doodle_left_alpha[64][74] = 1'b1; \
	doodle_left_alpha[64][75] = 1'b1; \
	doodle_left_alpha[64][76] = 1'b1; \
	doodle_left_alpha[64][77] = 1'b1; \
	doodle_left_alpha[64][78] = 1'b1; \
	doodle_left_alpha[64][79] = 1'b1; \
	doodle_left_alpha[65][0] = 1'b1; \
	doodle_left_alpha[65][1] = 1'b1; \
	doodle_left_alpha[65][2] = 1'b1; \
	doodle_left_alpha[65][3] = 1'b1; \
	doodle_left_alpha[65][4] = 1'b1; \
	doodle_left_alpha[65][5] = 1'b1; \
	doodle_left_alpha[65][6] = 1'b1; \
	doodle_left_alpha[65][7] = 1'b1; \
	doodle_left_alpha[65][8] = 1'b1; \
	doodle_left_alpha[65][9] = 1'b1; \
	doodle_left_alpha[65][10] = 1'b1; \
	doodle_left_alpha[65][11] = 1'b1; \
	doodle_left_alpha[65][12] = 1'b1; \
	doodle_left_alpha[65][13] = 1'b1; \
	doodle_left_alpha[65][14] = 1'b1; \
	doodle_left_alpha[65][15] = 1'b1; \
	doodle_left_alpha[65][16] = 1'b1; \
	doodle_left_alpha[65][17] = 1'b1; \
	doodle_left_alpha[65][18] = 1'b1; \
	doodle_left_alpha[65][19] = 1'b1; \
	doodle_left_alpha[65][20] = 1'b1; \
	doodle_left_alpha[65][21] = 1'b1; \
	doodle_left_alpha[65][22] = 1'b1; \
	doodle_left_alpha[65][23] = 1'b0; \
	doodle_left_alpha[65][24] = 1'b0; \
	doodle_left_alpha[65][25] = 1'b0; \
	doodle_left_alpha[65][26] = 1'b0; \
	doodle_left_alpha[65][27] = 1'b0; \
	doodle_left_alpha[65][28] = 1'b0; \
	doodle_left_alpha[65][29] = 1'b0; \
	doodle_left_alpha[65][30] = 1'b0; \
	doodle_left_alpha[65][31] = 1'b0; \
	doodle_left_alpha[65][32] = 1'b0; \
	doodle_left_alpha[65][33] = 1'b0; \
	doodle_left_alpha[65][34] = 1'b0; \
	doodle_left_alpha[65][35] = 1'b0; \
	doodle_left_alpha[65][36] = 1'b0; \
	doodle_left_alpha[65][37] = 1'b0; \
	doodle_left_alpha[65][38] = 1'b0; \
	doodle_left_alpha[65][39] = 1'b0; \
	doodle_left_alpha[65][40] = 1'b0; \
	doodle_left_alpha[65][41] = 1'b0; \
	doodle_left_alpha[65][42] = 1'b0; \
	doodle_left_alpha[65][43] = 1'b0; \
	doodle_left_alpha[65][44] = 1'b0; \
	doodle_left_alpha[65][45] = 1'b0; \
	doodle_left_alpha[65][46] = 1'b0; \
	doodle_left_alpha[65][47] = 1'b0; \
	doodle_left_alpha[65][48] = 1'b0; \
	doodle_left_alpha[65][49] = 1'b0; \
	doodle_left_alpha[65][50] = 1'b0; \
	doodle_left_alpha[65][51] = 1'b0; \
	doodle_left_alpha[65][52] = 1'b0; \
	doodle_left_alpha[65][53] = 1'b0; \
	doodle_left_alpha[65][54] = 1'b0; \
	doodle_left_alpha[65][55] = 1'b0; \
	doodle_left_alpha[65][56] = 1'b0; \
	doodle_left_alpha[65][57] = 1'b0; \
	doodle_left_alpha[65][58] = 1'b0; \
	doodle_left_alpha[65][59] = 1'b0; \
	doodle_left_alpha[65][60] = 1'b0; \
	doodle_left_alpha[65][61] = 1'b0; \
	doodle_left_alpha[65][62] = 1'b0; \
	doodle_left_alpha[65][63] = 1'b0; \
	doodle_left_alpha[65][64] = 1'b0; \
	doodle_left_alpha[65][65] = 1'b1; \
	doodle_left_alpha[65][66] = 1'b1; \
	doodle_left_alpha[65][67] = 1'b1; \
	doodle_left_alpha[65][68] = 1'b1; \
	doodle_left_alpha[65][69] = 1'b1; \
	doodle_left_alpha[65][70] = 1'b1; \
	doodle_left_alpha[65][71] = 1'b1; \
	doodle_left_alpha[65][72] = 1'b1; \
	doodle_left_alpha[65][73] = 1'b1; \
	doodle_left_alpha[65][74] = 1'b1; \
	doodle_left_alpha[65][75] = 1'b1; \
	doodle_left_alpha[65][76] = 1'b1; \
	doodle_left_alpha[65][77] = 1'b1; \
	doodle_left_alpha[65][78] = 1'b1; \
	doodle_left_alpha[65][79] = 1'b1; \
	doodle_left_alpha[66][0] = 1'b1; \
	doodle_left_alpha[66][1] = 1'b1; \
	doodle_left_alpha[66][2] = 1'b1; \
	doodle_left_alpha[66][3] = 1'b1; \
	doodle_left_alpha[66][4] = 1'b1; \
	doodle_left_alpha[66][5] = 1'b1; \
	doodle_left_alpha[66][6] = 1'b1; \
	doodle_left_alpha[66][7] = 1'b1; \
	doodle_left_alpha[66][8] = 1'b1; \
	doodle_left_alpha[66][9] = 1'b1; \
	doodle_left_alpha[66][10] = 1'b1; \
	doodle_left_alpha[66][11] = 1'b1; \
	doodle_left_alpha[66][12] = 1'b1; \
	doodle_left_alpha[66][13] = 1'b1; \
	doodle_left_alpha[66][14] = 1'b1; \
	doodle_left_alpha[66][15] = 1'b1; \
	doodle_left_alpha[66][16] = 1'b1; \
	doodle_left_alpha[66][17] = 1'b1; \
	doodle_left_alpha[66][18] = 1'b1; \
	doodle_left_alpha[66][19] = 1'b1; \
	doodle_left_alpha[66][20] = 1'b1; \
	doodle_left_alpha[66][21] = 1'b1; \
	doodle_left_alpha[66][22] = 1'b1; \
	doodle_left_alpha[66][23] = 1'b0; \
	doodle_left_alpha[66][24] = 1'b0; \
	doodle_left_alpha[66][25] = 1'b0; \
	doodle_left_alpha[66][26] = 1'b0; \
	doodle_left_alpha[66][27] = 1'b0; \
	doodle_left_alpha[66][28] = 1'b0; \
	doodle_left_alpha[66][29] = 1'b0; \
	doodle_left_alpha[66][30] = 1'b0; \
	doodle_left_alpha[66][31] = 1'b0; \
	doodle_left_alpha[66][32] = 1'b0; \
	doodle_left_alpha[66][33] = 1'b0; \
	doodle_left_alpha[66][34] = 1'b0; \
	doodle_left_alpha[66][35] = 1'b0; \
	doodle_left_alpha[66][36] = 1'b0; \
	doodle_left_alpha[66][37] = 1'b0; \
	doodle_left_alpha[66][38] = 1'b0; \
	doodle_left_alpha[66][39] = 1'b0; \
	doodle_left_alpha[66][40] = 1'b0; \
	doodle_left_alpha[66][41] = 1'b0; \
	doodle_left_alpha[66][42] = 1'b0; \
	doodle_left_alpha[66][43] = 1'b0; \
	doodle_left_alpha[66][44] = 1'b0; \
	doodle_left_alpha[66][45] = 1'b0; \
	doodle_left_alpha[66][46] = 1'b0; \
	doodle_left_alpha[66][47] = 1'b0; \
	doodle_left_alpha[66][48] = 1'b0; \
	doodle_left_alpha[66][49] = 1'b0; \
	doodle_left_alpha[66][50] = 1'b0; \
	doodle_left_alpha[66][51] = 1'b0; \
	doodle_left_alpha[66][52] = 1'b0; \
	doodle_left_alpha[66][53] = 1'b0; \
	doodle_left_alpha[66][54] = 1'b0; \
	doodle_left_alpha[66][55] = 1'b0; \
	doodle_left_alpha[66][56] = 1'b0; \
	doodle_left_alpha[66][57] = 1'b0; \
	doodle_left_alpha[66][58] = 1'b0; \
	doodle_left_alpha[66][59] = 1'b0; \
	doodle_left_alpha[66][60] = 1'b0; \
	doodle_left_alpha[66][61] = 1'b0; \
	doodle_left_alpha[66][62] = 1'b0; \
	doodle_left_alpha[66][63] = 1'b0; \
	doodle_left_alpha[66][64] = 1'b0; \
	doodle_left_alpha[66][65] = 1'b1; \
	doodle_left_alpha[66][66] = 1'b1; \
	doodle_left_alpha[66][67] = 1'b1; \
	doodle_left_alpha[66][68] = 1'b1; \
	doodle_left_alpha[66][69] = 1'b1; \
	doodle_left_alpha[66][70] = 1'b1; \
	doodle_left_alpha[66][71] = 1'b1; \
	doodle_left_alpha[66][72] = 1'b1; \
	doodle_left_alpha[66][73] = 1'b1; \
	doodle_left_alpha[66][74] = 1'b1; \
	doodle_left_alpha[66][75] = 1'b1; \
	doodle_left_alpha[66][76] = 1'b1; \
	doodle_left_alpha[66][77] = 1'b1; \
	doodle_left_alpha[66][78] = 1'b1; \
	doodle_left_alpha[66][79] = 1'b1; \
	doodle_left_alpha[67][0] = 1'b1; \
	doodle_left_alpha[67][1] = 1'b1; \
	doodle_left_alpha[67][2] = 1'b1; \
	doodle_left_alpha[67][3] = 1'b1; \
	doodle_left_alpha[67][4] = 1'b1; \
	doodle_left_alpha[67][5] = 1'b1; \
	doodle_left_alpha[67][6] = 1'b1; \
	doodle_left_alpha[67][7] = 1'b1; \
	doodle_left_alpha[67][8] = 1'b1; \
	doodle_left_alpha[67][9] = 1'b1; \
	doodle_left_alpha[67][10] = 1'b1; \
	doodle_left_alpha[67][11] = 1'b1; \
	doodle_left_alpha[67][12] = 1'b1; \
	doodle_left_alpha[67][13] = 1'b1; \
	doodle_left_alpha[67][14] = 1'b1; \
	doodle_left_alpha[67][15] = 1'b1; \
	doodle_left_alpha[67][16] = 1'b1; \
	doodle_left_alpha[67][17] = 1'b1; \
	doodle_left_alpha[67][18] = 1'b1; \
	doodle_left_alpha[67][19] = 1'b1; \
	doodle_left_alpha[67][20] = 1'b1; \
	doodle_left_alpha[67][21] = 1'b1; \
	doodle_left_alpha[67][22] = 1'b1; \
	doodle_left_alpha[67][23] = 1'b0; \
	doodle_left_alpha[67][24] = 1'b0; \
	doodle_left_alpha[67][25] = 1'b0; \
	doodle_left_alpha[67][26] = 1'b0; \
	doodle_left_alpha[67][27] = 1'b0; \
	doodle_left_alpha[67][28] = 1'b0; \
	doodle_left_alpha[67][29] = 1'b0; \
	doodle_left_alpha[67][30] = 1'b0; \
	doodle_left_alpha[67][31] = 1'b0; \
	doodle_left_alpha[67][32] = 1'b0; \
	doodle_left_alpha[67][33] = 1'b0; \
	doodle_left_alpha[67][34] = 1'b0; \
	doodle_left_alpha[67][35] = 1'b0; \
	doodle_left_alpha[67][36] = 1'b0; \
	doodle_left_alpha[67][37] = 1'b0; \
	doodle_left_alpha[67][38] = 1'b0; \
	doodle_left_alpha[67][39] = 1'b0; \
	doodle_left_alpha[67][40] = 1'b0; \
	doodle_left_alpha[67][41] = 1'b0; \
	doodle_left_alpha[67][42] = 1'b0; \
	doodle_left_alpha[67][43] = 1'b0; \
	doodle_left_alpha[67][44] = 1'b0; \
	doodle_left_alpha[67][45] = 1'b0; \
	doodle_left_alpha[67][46] = 1'b0; \
	doodle_left_alpha[67][47] = 1'b0; \
	doodle_left_alpha[67][48] = 1'b0; \
	doodle_left_alpha[67][49] = 1'b0; \
	doodle_left_alpha[67][50] = 1'b0; \
	doodle_left_alpha[67][51] = 1'b0; \
	doodle_left_alpha[67][52] = 1'b0; \
	doodle_left_alpha[67][53] = 1'b0; \
	doodle_left_alpha[67][54] = 1'b0; \
	doodle_left_alpha[67][55] = 1'b0; \
	doodle_left_alpha[67][56] = 1'b0; \
	doodle_left_alpha[67][57] = 1'b0; \
	doodle_left_alpha[67][58] = 1'b0; \
	doodle_left_alpha[67][59] = 1'b0; \
	doodle_left_alpha[67][60] = 1'b0; \
	doodle_left_alpha[67][61] = 1'b0; \
	doodle_left_alpha[67][62] = 1'b0; \
	doodle_left_alpha[67][63] = 1'b0; \
	doodle_left_alpha[67][64] = 1'b0; \
	doodle_left_alpha[67][65] = 1'b1; \
	doodle_left_alpha[67][66] = 1'b1; \
	doodle_left_alpha[67][67] = 1'b1; \
	doodle_left_alpha[67][68] = 1'b1; \
	doodle_left_alpha[67][69] = 1'b1; \
	doodle_left_alpha[67][70] = 1'b1; \
	doodle_left_alpha[67][71] = 1'b1; \
	doodle_left_alpha[67][72] = 1'b1; \
	doodle_left_alpha[67][73] = 1'b1; \
	doodle_left_alpha[67][74] = 1'b1; \
	doodle_left_alpha[67][75] = 1'b1; \
	doodle_left_alpha[67][76] = 1'b1; \
	doodle_left_alpha[67][77] = 1'b1; \
	doodle_left_alpha[67][78] = 1'b1; \
	doodle_left_alpha[67][79] = 1'b1; \
	doodle_left_alpha[68][0] = 1'b1; \
	doodle_left_alpha[68][1] = 1'b1; \
	doodle_left_alpha[68][2] = 1'b1; \
	doodle_left_alpha[68][3] = 1'b1; \
	doodle_left_alpha[68][4] = 1'b1; \
	doodle_left_alpha[68][5] = 1'b1; \
	doodle_left_alpha[68][6] = 1'b1; \
	doodle_left_alpha[68][7] = 1'b1; \
	doodle_left_alpha[68][8] = 1'b1; \
	doodle_left_alpha[68][9] = 1'b1; \
	doodle_left_alpha[68][10] = 1'b1; \
	doodle_left_alpha[68][11] = 1'b1; \
	doodle_left_alpha[68][12] = 1'b1; \
	doodle_left_alpha[68][13] = 1'b1; \
	doodle_left_alpha[68][14] = 1'b1; \
	doodle_left_alpha[68][15] = 1'b1; \
	doodle_left_alpha[68][16] = 1'b1; \
	doodle_left_alpha[68][17] = 1'b1; \
	doodle_left_alpha[68][18] = 1'b1; \
	doodle_left_alpha[68][19] = 1'b1; \
	doodle_left_alpha[68][20] = 1'b1; \
	doodle_left_alpha[68][21] = 1'b1; \
	doodle_left_alpha[68][22] = 1'b1; \
	doodle_left_alpha[68][23] = 1'b1; \
	doodle_left_alpha[68][24] = 1'b1; \
	doodle_left_alpha[68][25] = 1'b1; \
	doodle_left_alpha[68][26] = 1'b1; \
	doodle_left_alpha[68][27] = 1'b0; \
	doodle_left_alpha[68][28] = 1'b0; \
	doodle_left_alpha[68][29] = 1'b0; \
	doodle_left_alpha[68][30] = 1'b0; \
	doodle_left_alpha[68][31] = 1'b1; \
	doodle_left_alpha[68][32] = 1'b1; \
	doodle_left_alpha[68][33] = 1'b1; \
	doodle_left_alpha[68][34] = 1'b1; \
	doodle_left_alpha[68][35] = 1'b1; \
	doodle_left_alpha[68][36] = 1'b1; \
	doodle_left_alpha[68][37] = 1'b0; \
	doodle_left_alpha[68][38] = 1'b0; \
	doodle_left_alpha[68][39] = 1'b0; \
	doodle_left_alpha[68][40] = 1'b0; \
	doodle_left_alpha[68][41] = 1'b1; \
	doodle_left_alpha[68][42] = 1'b1; \
	doodle_left_alpha[68][43] = 1'b1; \
	doodle_left_alpha[68][44] = 1'b1; \
	doodle_left_alpha[68][45] = 1'b1; \
	doodle_left_alpha[68][46] = 1'b1; \
	doodle_left_alpha[68][47] = 1'b0; \
	doodle_left_alpha[68][48] = 1'b0; \
	doodle_left_alpha[68][49] = 1'b0; \
	doodle_left_alpha[68][50] = 1'b0; \
	doodle_left_alpha[68][51] = 1'b1; \
	doodle_left_alpha[68][52] = 1'b1; \
	doodle_left_alpha[68][53] = 1'b1; \
	doodle_left_alpha[68][54] = 1'b1; \
	doodle_left_alpha[68][55] = 1'b1; \
	doodle_left_alpha[68][56] = 1'b1; \
	doodle_left_alpha[68][57] = 1'b0; \
	doodle_left_alpha[68][58] = 1'b0; \
	doodle_left_alpha[68][59] = 1'b0; \
	doodle_left_alpha[68][60] = 1'b0; \
	doodle_left_alpha[68][61] = 1'b1; \
	doodle_left_alpha[68][62] = 1'b1; \
	doodle_left_alpha[68][63] = 1'b1; \
	doodle_left_alpha[68][64] = 1'b1; \
	doodle_left_alpha[68][65] = 1'b1; \
	doodle_left_alpha[68][66] = 1'b1; \
	doodle_left_alpha[68][67] = 1'b1; \
	doodle_left_alpha[68][68] = 1'b1; \
	doodle_left_alpha[68][69] = 1'b1; \
	doodle_left_alpha[68][70] = 1'b1; \
	doodle_left_alpha[68][71] = 1'b1; \
	doodle_left_alpha[68][72] = 1'b1; \
	doodle_left_alpha[68][73] = 1'b1; \
	doodle_left_alpha[68][74] = 1'b1; \
	doodle_left_alpha[68][75] = 1'b1; \
	doodle_left_alpha[68][76] = 1'b1; \
	doodle_left_alpha[68][77] = 1'b1; \
	doodle_left_alpha[68][78] = 1'b1; \
	doodle_left_alpha[68][79] = 1'b1; \
	doodle_left_alpha[69][0] = 1'b1; \
	doodle_left_alpha[69][1] = 1'b1; \
	doodle_left_alpha[69][2] = 1'b1; \
	doodle_left_alpha[69][3] = 1'b1; \
	doodle_left_alpha[69][4] = 1'b1; \
	doodle_left_alpha[69][5] = 1'b1; \
	doodle_left_alpha[69][6] = 1'b1; \
	doodle_left_alpha[69][7] = 1'b1; \
	doodle_left_alpha[69][8] = 1'b1; \
	doodle_left_alpha[69][9] = 1'b1; \
	doodle_left_alpha[69][10] = 1'b1; \
	doodle_left_alpha[69][11] = 1'b1; \
	doodle_left_alpha[69][12] = 1'b1; \
	doodle_left_alpha[69][13] = 1'b1; \
	doodle_left_alpha[69][14] = 1'b1; \
	doodle_left_alpha[69][15] = 1'b1; \
	doodle_left_alpha[69][16] = 1'b1; \
	doodle_left_alpha[69][17] = 1'b1; \
	doodle_left_alpha[69][18] = 1'b1; \
	doodle_left_alpha[69][19] = 1'b1; \
	doodle_left_alpha[69][20] = 1'b1; \
	doodle_left_alpha[69][21] = 1'b1; \
	doodle_left_alpha[69][22] = 1'b1; \
	doodle_left_alpha[69][23] = 1'b1; \
	doodle_left_alpha[69][24] = 1'b1; \
	doodle_left_alpha[69][25] = 1'b1; \
	doodle_left_alpha[69][26] = 1'b1; \
	doodle_left_alpha[69][27] = 1'b0; \
	doodle_left_alpha[69][28] = 1'b0; \
	doodle_left_alpha[69][29] = 1'b0; \
	doodle_left_alpha[69][30] = 1'b0; \
	doodle_left_alpha[69][31] = 1'b1; \
	doodle_left_alpha[69][32] = 1'b1; \
	doodle_left_alpha[69][33] = 1'b1; \
	doodle_left_alpha[69][34] = 1'b1; \
	doodle_left_alpha[69][35] = 1'b1; \
	doodle_left_alpha[69][36] = 1'b1; \
	doodle_left_alpha[69][37] = 1'b0; \
	doodle_left_alpha[69][38] = 1'b0; \
	doodle_left_alpha[69][39] = 1'b0; \
	doodle_left_alpha[69][40] = 1'b0; \
	doodle_left_alpha[69][41] = 1'b1; \
	doodle_left_alpha[69][42] = 1'b1; \
	doodle_left_alpha[69][43] = 1'b1; \
	doodle_left_alpha[69][44] = 1'b1; \
	doodle_left_alpha[69][45] = 1'b1; \
	doodle_left_alpha[69][46] = 1'b1; \
	doodle_left_alpha[69][47] = 1'b0; \
	doodle_left_alpha[69][48] = 1'b0; \
	doodle_left_alpha[69][49] = 1'b0; \
	doodle_left_alpha[69][50] = 1'b0; \
	doodle_left_alpha[69][51] = 1'b1; \
	doodle_left_alpha[69][52] = 1'b1; \
	doodle_left_alpha[69][53] = 1'b1; \
	doodle_left_alpha[69][54] = 1'b1; \
	doodle_left_alpha[69][55] = 1'b1; \
	doodle_left_alpha[69][56] = 1'b1; \
	doodle_left_alpha[69][57] = 1'b0; \
	doodle_left_alpha[69][58] = 1'b0; \
	doodle_left_alpha[69][59] = 1'b0; \
	doodle_left_alpha[69][60] = 1'b0; \
	doodle_left_alpha[69][61] = 1'b1; \
	doodle_left_alpha[69][62] = 1'b1; \
	doodle_left_alpha[69][63] = 1'b1; \
	doodle_left_alpha[69][64] = 1'b1; \
	doodle_left_alpha[69][65] = 1'b1; \
	doodle_left_alpha[69][66] = 1'b1; \
	doodle_left_alpha[69][67] = 1'b1; \
	doodle_left_alpha[69][68] = 1'b1; \
	doodle_left_alpha[69][69] = 1'b1; \
	doodle_left_alpha[69][70] = 1'b1; \
	doodle_left_alpha[69][71] = 1'b1; \
	doodle_left_alpha[69][72] = 1'b1; \
	doodle_left_alpha[69][73] = 1'b1; \
	doodle_left_alpha[69][74] = 1'b1; \
	doodle_left_alpha[69][75] = 1'b1; \
	doodle_left_alpha[69][76] = 1'b1; \
	doodle_left_alpha[69][77] = 1'b1; \
	doodle_left_alpha[69][78] = 1'b1; \
	doodle_left_alpha[69][79] = 1'b1; \
	doodle_left_alpha[70][0] = 1'b1; \
	doodle_left_alpha[70][1] = 1'b1; \
	doodle_left_alpha[70][2] = 1'b1; \
	doodle_left_alpha[70][3] = 1'b1; \
	doodle_left_alpha[70][4] = 1'b1; \
	doodle_left_alpha[70][5] = 1'b1; \
	doodle_left_alpha[70][6] = 1'b1; \
	doodle_left_alpha[70][7] = 1'b1; \
	doodle_left_alpha[70][8] = 1'b1; \
	doodle_left_alpha[70][9] = 1'b1; \
	doodle_left_alpha[70][10] = 1'b1; \
	doodle_left_alpha[70][11] = 1'b1; \
	doodle_left_alpha[70][12] = 1'b1; \
	doodle_left_alpha[70][13] = 1'b1; \
	doodle_left_alpha[70][14] = 1'b1; \
	doodle_left_alpha[70][15] = 1'b1; \
	doodle_left_alpha[70][16] = 1'b1; \
	doodle_left_alpha[70][17] = 1'b1; \
	doodle_left_alpha[70][18] = 1'b1; \
	doodle_left_alpha[70][19] = 1'b1; \
	doodle_left_alpha[70][20] = 1'b1; \
	doodle_left_alpha[70][21] = 1'b1; \
	doodle_left_alpha[70][22] = 1'b1; \
	doodle_left_alpha[70][23] = 1'b1; \
	doodle_left_alpha[70][24] = 1'b1; \
	doodle_left_alpha[70][25] = 1'b1; \
	doodle_left_alpha[70][26] = 1'b1; \
	doodle_left_alpha[70][27] = 1'b0; \
	doodle_left_alpha[70][28] = 1'b0; \
	doodle_left_alpha[70][29] = 1'b0; \
	doodle_left_alpha[70][30] = 1'b0; \
	doodle_left_alpha[70][31] = 1'b1; \
	doodle_left_alpha[70][32] = 1'b1; \
	doodle_left_alpha[70][33] = 1'b1; \
	doodle_left_alpha[70][34] = 1'b1; \
	doodle_left_alpha[70][35] = 1'b1; \
	doodle_left_alpha[70][36] = 1'b1; \
	doodle_left_alpha[70][37] = 1'b0; \
	doodle_left_alpha[70][38] = 1'b0; \
	doodle_left_alpha[70][39] = 1'b0; \
	doodle_left_alpha[70][40] = 1'b0; \
	doodle_left_alpha[70][41] = 1'b1; \
	doodle_left_alpha[70][42] = 1'b1; \
	doodle_left_alpha[70][43] = 1'b1; \
	doodle_left_alpha[70][44] = 1'b1; \
	doodle_left_alpha[70][45] = 1'b1; \
	doodle_left_alpha[70][46] = 1'b1; \
	doodle_left_alpha[70][47] = 1'b0; \
	doodle_left_alpha[70][48] = 1'b0; \
	doodle_left_alpha[70][49] = 1'b0; \
	doodle_left_alpha[70][50] = 1'b0; \
	doodle_left_alpha[70][51] = 1'b1; \
	doodle_left_alpha[70][52] = 1'b1; \
	doodle_left_alpha[70][53] = 1'b1; \
	doodle_left_alpha[70][54] = 1'b1; \
	doodle_left_alpha[70][55] = 1'b1; \
	doodle_left_alpha[70][56] = 1'b1; \
	doodle_left_alpha[70][57] = 1'b0; \
	doodle_left_alpha[70][58] = 1'b0; \
	doodle_left_alpha[70][59] = 1'b0; \
	doodle_left_alpha[70][60] = 1'b0; \
	doodle_left_alpha[70][61] = 1'b1; \
	doodle_left_alpha[70][62] = 1'b1; \
	doodle_left_alpha[70][63] = 1'b1; \
	doodle_left_alpha[70][64] = 1'b1; \
	doodle_left_alpha[70][65] = 1'b1; \
	doodle_left_alpha[70][66] = 1'b1; \
	doodle_left_alpha[70][67] = 1'b1; \
	doodle_left_alpha[70][68] = 1'b1; \
	doodle_left_alpha[70][69] = 1'b1; \
	doodle_left_alpha[70][70] = 1'b1; \
	doodle_left_alpha[70][71] = 1'b1; \
	doodle_left_alpha[70][72] = 1'b1; \
	doodle_left_alpha[70][73] = 1'b1; \
	doodle_left_alpha[70][74] = 1'b1; \
	doodle_left_alpha[70][75] = 1'b1; \
	doodle_left_alpha[70][76] = 1'b1; \
	doodle_left_alpha[70][77] = 1'b1; \
	doodle_left_alpha[70][78] = 1'b1; \
	doodle_left_alpha[70][79] = 1'b1; \
	doodle_left_alpha[71][0] = 1'b1; \
	doodle_left_alpha[71][1] = 1'b1; \
	doodle_left_alpha[71][2] = 1'b1; \
	doodle_left_alpha[71][3] = 1'b1; \
	doodle_left_alpha[71][4] = 1'b1; \
	doodle_left_alpha[71][5] = 1'b1; \
	doodle_left_alpha[71][6] = 1'b1; \
	doodle_left_alpha[71][7] = 1'b1; \
	doodle_left_alpha[71][8] = 1'b1; \
	doodle_left_alpha[71][9] = 1'b1; \
	doodle_left_alpha[71][10] = 1'b1; \
	doodle_left_alpha[71][11] = 1'b1; \
	doodle_left_alpha[71][12] = 1'b1; \
	doodle_left_alpha[71][13] = 1'b1; \
	doodle_left_alpha[71][14] = 1'b1; \
	doodle_left_alpha[71][15] = 1'b1; \
	doodle_left_alpha[71][16] = 1'b1; \
	doodle_left_alpha[71][17] = 1'b1; \
	doodle_left_alpha[71][18] = 1'b1; \
	doodle_left_alpha[71][19] = 1'b1; \
	doodle_left_alpha[71][20] = 1'b1; \
	doodle_left_alpha[71][21] = 1'b1; \
	doodle_left_alpha[71][22] = 1'b1; \
	doodle_left_alpha[71][23] = 1'b1; \
	doodle_left_alpha[71][24] = 1'b1; \
	doodle_left_alpha[71][25] = 1'b1; \
	doodle_left_alpha[71][26] = 1'b1; \
	doodle_left_alpha[71][27] = 1'b0; \
	doodle_left_alpha[71][28] = 1'b0; \
	doodle_left_alpha[71][29] = 1'b0; \
	doodle_left_alpha[71][30] = 1'b0; \
	doodle_left_alpha[71][31] = 1'b1; \
	doodle_left_alpha[71][32] = 1'b1; \
	doodle_left_alpha[71][33] = 1'b1; \
	doodle_left_alpha[71][34] = 1'b1; \
	doodle_left_alpha[71][35] = 1'b1; \
	doodle_left_alpha[71][36] = 1'b1; \
	doodle_left_alpha[71][37] = 1'b0; \
	doodle_left_alpha[71][38] = 1'b0; \
	doodle_left_alpha[71][39] = 1'b0; \
	doodle_left_alpha[71][40] = 1'b0; \
	doodle_left_alpha[71][41] = 1'b1; \
	doodle_left_alpha[71][42] = 1'b1; \
	doodle_left_alpha[71][43] = 1'b1; \
	doodle_left_alpha[71][44] = 1'b1; \
	doodle_left_alpha[71][45] = 1'b1; \
	doodle_left_alpha[71][46] = 1'b1; \
	doodle_left_alpha[71][47] = 1'b0; \
	doodle_left_alpha[71][48] = 1'b0; \
	doodle_left_alpha[71][49] = 1'b0; \
	doodle_left_alpha[71][50] = 1'b0; \
	doodle_left_alpha[71][51] = 1'b1; \
	doodle_left_alpha[71][52] = 1'b1; \
	doodle_left_alpha[71][53] = 1'b1; \
	doodle_left_alpha[71][54] = 1'b1; \
	doodle_left_alpha[71][55] = 1'b1; \
	doodle_left_alpha[71][56] = 1'b1; \
	doodle_left_alpha[71][57] = 1'b0; \
	doodle_left_alpha[71][58] = 1'b0; \
	doodle_left_alpha[71][59] = 1'b0; \
	doodle_left_alpha[71][60] = 1'b0; \
	doodle_left_alpha[71][61] = 1'b1; \
	doodle_left_alpha[71][62] = 1'b1; \
	doodle_left_alpha[71][63] = 1'b1; \
	doodle_left_alpha[71][64] = 1'b1; \
	doodle_left_alpha[71][65] = 1'b1; \
	doodle_left_alpha[71][66] = 1'b1; \
	doodle_left_alpha[71][67] = 1'b1; \
	doodle_left_alpha[71][68] = 1'b1; \
	doodle_left_alpha[71][69] = 1'b1; \
	doodle_left_alpha[71][70] = 1'b1; \
	doodle_left_alpha[71][71] = 1'b1; \
	doodle_left_alpha[71][72] = 1'b1; \
	doodle_left_alpha[71][73] = 1'b1; \
	doodle_left_alpha[71][74] = 1'b1; \
	doodle_left_alpha[71][75] = 1'b1; \
	doodle_left_alpha[71][76] = 1'b1; \
	doodle_left_alpha[71][77] = 1'b1; \
	doodle_left_alpha[71][78] = 1'b1; \
	doodle_left_alpha[71][79] = 1'b1; \
	doodle_left_alpha[72][0] = 1'b1; \
	doodle_left_alpha[72][1] = 1'b1; \
	doodle_left_alpha[72][2] = 1'b1; \
	doodle_left_alpha[72][3] = 1'b1; \
	doodle_left_alpha[72][4] = 1'b1; \
	doodle_left_alpha[72][5] = 1'b1; \
	doodle_left_alpha[72][6] = 1'b1; \
	doodle_left_alpha[72][7] = 1'b1; \
	doodle_left_alpha[72][8] = 1'b1; \
	doodle_left_alpha[72][9] = 1'b1; \
	doodle_left_alpha[72][10] = 1'b1; \
	doodle_left_alpha[72][11] = 1'b1; \
	doodle_left_alpha[72][12] = 1'b1; \
	doodle_left_alpha[72][13] = 1'b1; \
	doodle_left_alpha[72][14] = 1'b1; \
	doodle_left_alpha[72][15] = 1'b1; \
	doodle_left_alpha[72][16] = 1'b1; \
	doodle_left_alpha[72][17] = 1'b1; \
	doodle_left_alpha[72][18] = 1'b1; \
	doodle_left_alpha[72][19] = 1'b1; \
	doodle_left_alpha[72][20] = 1'b1; \
	doodle_left_alpha[72][21] = 1'b1; \
	doodle_left_alpha[72][22] = 1'b1; \
	doodle_left_alpha[72][23] = 1'b1; \
	doodle_left_alpha[72][24] = 1'b1; \
	doodle_left_alpha[72][25] = 1'b1; \
	doodle_left_alpha[72][26] = 1'b1; \
	doodle_left_alpha[72][27] = 1'b0; \
	doodle_left_alpha[72][28] = 1'b0; \
	doodle_left_alpha[72][29] = 1'b0; \
	doodle_left_alpha[72][30] = 1'b0; \
	doodle_left_alpha[72][31] = 1'b1; \
	doodle_left_alpha[72][32] = 1'b1; \
	doodle_left_alpha[72][33] = 1'b1; \
	doodle_left_alpha[72][34] = 1'b1; \
	doodle_left_alpha[72][35] = 1'b1; \
	doodle_left_alpha[72][36] = 1'b1; \
	doodle_left_alpha[72][37] = 1'b0; \
	doodle_left_alpha[72][38] = 1'b0; \
	doodle_left_alpha[72][39] = 1'b0; \
	doodle_left_alpha[72][40] = 1'b0; \
	doodle_left_alpha[72][41] = 1'b1; \
	doodle_left_alpha[72][42] = 1'b1; \
	doodle_left_alpha[72][43] = 1'b1; \
	doodle_left_alpha[72][44] = 1'b1; \
	doodle_left_alpha[72][45] = 1'b1; \
	doodle_left_alpha[72][46] = 1'b1; \
	doodle_left_alpha[72][47] = 1'b0; \
	doodle_left_alpha[72][48] = 1'b0; \
	doodle_left_alpha[72][49] = 1'b0; \
	doodle_left_alpha[72][50] = 1'b0; \
	doodle_left_alpha[72][51] = 1'b1; \
	doodle_left_alpha[72][52] = 1'b1; \
	doodle_left_alpha[72][53] = 1'b1; \
	doodle_left_alpha[72][54] = 1'b1; \
	doodle_left_alpha[72][55] = 1'b1; \
	doodle_left_alpha[72][56] = 1'b1; \
	doodle_left_alpha[72][57] = 1'b0; \
	doodle_left_alpha[72][58] = 1'b0; \
	doodle_left_alpha[72][59] = 1'b0; \
	doodle_left_alpha[72][60] = 1'b0; \
	doodle_left_alpha[72][61] = 1'b1; \
	doodle_left_alpha[72][62] = 1'b1; \
	doodle_left_alpha[72][63] = 1'b1; \
	doodle_left_alpha[72][64] = 1'b1; \
	doodle_left_alpha[72][65] = 1'b1; \
	doodle_left_alpha[72][66] = 1'b1; \
	doodle_left_alpha[72][67] = 1'b1; \
	doodle_left_alpha[72][68] = 1'b1; \
	doodle_left_alpha[72][69] = 1'b1; \
	doodle_left_alpha[72][70] = 1'b1; \
	doodle_left_alpha[72][71] = 1'b1; \
	doodle_left_alpha[72][72] = 1'b1; \
	doodle_left_alpha[72][73] = 1'b1; \
	doodle_left_alpha[72][74] = 1'b1; \
	doodle_left_alpha[72][75] = 1'b1; \
	doodle_left_alpha[72][76] = 1'b1; \
	doodle_left_alpha[72][77] = 1'b1; \
	doodle_left_alpha[72][78] = 1'b1; \
	doodle_left_alpha[72][79] = 1'b1; \
	doodle_left_alpha[73][0] = 1'b1; \
	doodle_left_alpha[73][1] = 1'b1; \
	doodle_left_alpha[73][2] = 1'b1; \
	doodle_left_alpha[73][3] = 1'b1; \
	doodle_left_alpha[73][4] = 1'b1; \
	doodle_left_alpha[73][5] = 1'b1; \
	doodle_left_alpha[73][6] = 1'b1; \
	doodle_left_alpha[73][7] = 1'b1; \
	doodle_left_alpha[73][8] = 1'b1; \
	doodle_left_alpha[73][9] = 1'b1; \
	doodle_left_alpha[73][10] = 1'b1; \
	doodle_left_alpha[73][11] = 1'b1; \
	doodle_left_alpha[73][12] = 1'b1; \
	doodle_left_alpha[73][13] = 1'b1; \
	doodle_left_alpha[73][14] = 1'b1; \
	doodle_left_alpha[73][15] = 1'b1; \
	doodle_left_alpha[73][16] = 1'b1; \
	doodle_left_alpha[73][17] = 1'b1; \
	doodle_left_alpha[73][18] = 1'b1; \
	doodle_left_alpha[73][19] = 1'b1; \
	doodle_left_alpha[73][20] = 1'b1; \
	doodle_left_alpha[73][21] = 1'b1; \
	doodle_left_alpha[73][22] = 1'b1; \
	doodle_left_alpha[73][23] = 1'b1; \
	doodle_left_alpha[73][24] = 1'b1; \
	doodle_left_alpha[73][25] = 1'b1; \
	doodle_left_alpha[73][26] = 1'b1; \
	doodle_left_alpha[73][27] = 1'b0; \
	doodle_left_alpha[73][28] = 1'b0; \
	doodle_left_alpha[73][29] = 1'b0; \
	doodle_left_alpha[73][30] = 1'b0; \
	doodle_left_alpha[73][31] = 1'b1; \
	doodle_left_alpha[73][32] = 1'b1; \
	doodle_left_alpha[73][33] = 1'b1; \
	doodle_left_alpha[73][34] = 1'b1; \
	doodle_left_alpha[73][35] = 1'b1; \
	doodle_left_alpha[73][36] = 1'b1; \
	doodle_left_alpha[73][37] = 1'b0; \
	doodle_left_alpha[73][38] = 1'b0; \
	doodle_left_alpha[73][39] = 1'b0; \
	doodle_left_alpha[73][40] = 1'b0; \
	doodle_left_alpha[73][41] = 1'b1; \
	doodle_left_alpha[73][42] = 1'b1; \
	doodle_left_alpha[73][43] = 1'b1; \
	doodle_left_alpha[73][44] = 1'b1; \
	doodle_left_alpha[73][45] = 1'b1; \
	doodle_left_alpha[73][46] = 1'b1; \
	doodle_left_alpha[73][47] = 1'b0; \
	doodle_left_alpha[73][48] = 1'b0; \
	doodle_left_alpha[73][49] = 1'b0; \
	doodle_left_alpha[73][50] = 1'b0; \
	doodle_left_alpha[73][51] = 1'b1; \
	doodle_left_alpha[73][52] = 1'b1; \
	doodle_left_alpha[73][53] = 1'b1; \
	doodle_left_alpha[73][54] = 1'b1; \
	doodle_left_alpha[73][55] = 1'b1; \
	doodle_left_alpha[73][56] = 1'b1; \
	doodle_left_alpha[73][57] = 1'b0; \
	doodle_left_alpha[73][58] = 1'b0; \
	doodle_left_alpha[73][59] = 1'b0; \
	doodle_left_alpha[73][60] = 1'b0; \
	doodle_left_alpha[73][61] = 1'b1; \
	doodle_left_alpha[73][62] = 1'b1; \
	doodle_left_alpha[73][63] = 1'b1; \
	doodle_left_alpha[73][64] = 1'b1; \
	doodle_left_alpha[73][65] = 1'b1; \
	doodle_left_alpha[73][66] = 1'b1; \
	doodle_left_alpha[73][67] = 1'b1; \
	doodle_left_alpha[73][68] = 1'b1; \
	doodle_left_alpha[73][69] = 1'b1; \
	doodle_left_alpha[73][70] = 1'b1; \
	doodle_left_alpha[73][71] = 1'b1; \
	doodle_left_alpha[73][72] = 1'b1; \
	doodle_left_alpha[73][73] = 1'b1; \
	doodle_left_alpha[73][74] = 1'b1; \
	doodle_left_alpha[73][75] = 1'b1; \
	doodle_left_alpha[73][76] = 1'b1; \
	doodle_left_alpha[73][77] = 1'b1; \
	doodle_left_alpha[73][78] = 1'b1; \
	doodle_left_alpha[73][79] = 1'b1; \
	doodle_left_alpha[74][0] = 1'b1; \
	doodle_left_alpha[74][1] = 1'b1; \
	doodle_left_alpha[74][2] = 1'b1; \
	doodle_left_alpha[74][3] = 1'b1; \
	doodle_left_alpha[74][4] = 1'b1; \
	doodle_left_alpha[74][5] = 1'b1; \
	doodle_left_alpha[74][6] = 1'b1; \
	doodle_left_alpha[74][7] = 1'b1; \
	doodle_left_alpha[74][8] = 1'b1; \
	doodle_left_alpha[74][9] = 1'b1; \
	doodle_left_alpha[74][10] = 1'b1; \
	doodle_left_alpha[74][11] = 1'b1; \
	doodle_left_alpha[74][12] = 1'b1; \
	doodle_left_alpha[74][13] = 1'b1; \
	doodle_left_alpha[74][14] = 1'b1; \
	doodle_left_alpha[74][15] = 1'b1; \
	doodle_left_alpha[74][16] = 1'b1; \
	doodle_left_alpha[74][17] = 1'b1; \
	doodle_left_alpha[74][18] = 1'b1; \
	doodle_left_alpha[74][19] = 1'b1; \
	doodle_left_alpha[74][20] = 1'b1; \
	doodle_left_alpha[74][21] = 1'b1; \
	doodle_left_alpha[74][22] = 1'b1; \
	doodle_left_alpha[74][23] = 1'b1; \
	doodle_left_alpha[74][24] = 1'b1; \
	doodle_left_alpha[74][25] = 1'b1; \
	doodle_left_alpha[74][26] = 1'b1; \
	doodle_left_alpha[74][27] = 1'b0; \
	doodle_left_alpha[74][28] = 1'b0; \
	doodle_left_alpha[74][29] = 1'b0; \
	doodle_left_alpha[74][30] = 1'b0; \
	doodle_left_alpha[74][31] = 1'b1; \
	doodle_left_alpha[74][32] = 1'b1; \
	doodle_left_alpha[74][33] = 1'b1; \
	doodle_left_alpha[74][34] = 1'b1; \
	doodle_left_alpha[74][35] = 1'b1; \
	doodle_left_alpha[74][36] = 1'b1; \
	doodle_left_alpha[74][37] = 1'b0; \
	doodle_left_alpha[74][38] = 1'b0; \
	doodle_left_alpha[74][39] = 1'b0; \
	doodle_left_alpha[74][40] = 1'b0; \
	doodle_left_alpha[74][41] = 1'b1; \
	doodle_left_alpha[74][42] = 1'b1; \
	doodle_left_alpha[74][43] = 1'b1; \
	doodle_left_alpha[74][44] = 1'b1; \
	doodle_left_alpha[74][45] = 1'b1; \
	doodle_left_alpha[74][46] = 1'b1; \
	doodle_left_alpha[74][47] = 1'b0; \
	doodle_left_alpha[74][48] = 1'b0; \
	doodle_left_alpha[74][49] = 1'b0; \
	doodle_left_alpha[74][50] = 1'b0; \
	doodle_left_alpha[74][51] = 1'b1; \
	doodle_left_alpha[74][52] = 1'b1; \
	doodle_left_alpha[74][53] = 1'b1; \
	doodle_left_alpha[74][54] = 1'b1; \
	doodle_left_alpha[74][55] = 1'b1; \
	doodle_left_alpha[74][56] = 1'b1; \
	doodle_left_alpha[74][57] = 1'b0; \
	doodle_left_alpha[74][58] = 1'b0; \
	doodle_left_alpha[74][59] = 1'b0; \
	doodle_left_alpha[74][60] = 1'b0; \
	doodle_left_alpha[74][61] = 1'b1; \
	doodle_left_alpha[74][62] = 1'b1; \
	doodle_left_alpha[74][63] = 1'b1; \
	doodle_left_alpha[74][64] = 1'b1; \
	doodle_left_alpha[74][65] = 1'b1; \
	doodle_left_alpha[74][66] = 1'b1; \
	doodle_left_alpha[74][67] = 1'b1; \
	doodle_left_alpha[74][68] = 1'b1; \
	doodle_left_alpha[74][69] = 1'b1; \
	doodle_left_alpha[74][70] = 1'b1; \
	doodle_left_alpha[74][71] = 1'b1; \
	doodle_left_alpha[74][72] = 1'b1; \
	doodle_left_alpha[74][73] = 1'b1; \
	doodle_left_alpha[74][74] = 1'b1; \
	doodle_left_alpha[74][75] = 1'b1; \
	doodle_left_alpha[74][76] = 1'b1; \
	doodle_left_alpha[74][77] = 1'b1; \
	doodle_left_alpha[74][78] = 1'b1; \
	doodle_left_alpha[74][79] = 1'b1; \
	doodle_left_alpha[75][0] = 1'b1; \
	doodle_left_alpha[75][1] = 1'b1; \
	doodle_left_alpha[75][2] = 1'b1; \
	doodle_left_alpha[75][3] = 1'b1; \
	doodle_left_alpha[75][4] = 1'b1; \
	doodle_left_alpha[75][5] = 1'b1; \
	doodle_left_alpha[75][6] = 1'b1; \
	doodle_left_alpha[75][7] = 1'b1; \
	doodle_left_alpha[75][8] = 1'b1; \
	doodle_left_alpha[75][9] = 1'b1; \
	doodle_left_alpha[75][10] = 1'b1; \
	doodle_left_alpha[75][11] = 1'b1; \
	doodle_left_alpha[75][12] = 1'b1; \
	doodle_left_alpha[75][13] = 1'b1; \
	doodle_left_alpha[75][14] = 1'b1; \
	doodle_left_alpha[75][15] = 1'b1; \
	doodle_left_alpha[75][16] = 1'b1; \
	doodle_left_alpha[75][17] = 1'b1; \
	doodle_left_alpha[75][18] = 1'b1; \
	doodle_left_alpha[75][19] = 1'b1; \
	doodle_left_alpha[75][20] = 1'b1; \
	doodle_left_alpha[75][21] = 1'b1; \
	doodle_left_alpha[75][22] = 1'b1; \
	doodle_left_alpha[75][23] = 1'b1; \
	doodle_left_alpha[75][24] = 1'b1; \
	doodle_left_alpha[75][25] = 1'b1; \
	doodle_left_alpha[75][26] = 1'b1; \
	doodle_left_alpha[75][27] = 1'b0; \
	doodle_left_alpha[75][28] = 1'b0; \
	doodle_left_alpha[75][29] = 1'b0; \
	doodle_left_alpha[75][30] = 1'b0; \
	doodle_left_alpha[75][31] = 1'b1; \
	doodle_left_alpha[75][32] = 1'b1; \
	doodle_left_alpha[75][33] = 1'b1; \
	doodle_left_alpha[75][34] = 1'b1; \
	doodle_left_alpha[75][35] = 1'b1; \
	doodle_left_alpha[75][36] = 1'b1; \
	doodle_left_alpha[75][37] = 1'b0; \
	doodle_left_alpha[75][38] = 1'b0; \
	doodle_left_alpha[75][39] = 1'b0; \
	doodle_left_alpha[75][40] = 1'b0; \
	doodle_left_alpha[75][41] = 1'b1; \
	doodle_left_alpha[75][42] = 1'b1; \
	doodle_left_alpha[75][43] = 1'b1; \
	doodle_left_alpha[75][44] = 1'b1; \
	doodle_left_alpha[75][45] = 1'b1; \
	doodle_left_alpha[75][46] = 1'b1; \
	doodle_left_alpha[75][47] = 1'b0; \
	doodle_left_alpha[75][48] = 1'b0; \
	doodle_left_alpha[75][49] = 1'b0; \
	doodle_left_alpha[75][50] = 1'b0; \
	doodle_left_alpha[75][51] = 1'b1; \
	doodle_left_alpha[75][52] = 1'b1; \
	doodle_left_alpha[75][53] = 1'b1; \
	doodle_left_alpha[75][54] = 1'b1; \
	doodle_left_alpha[75][55] = 1'b1; \
	doodle_left_alpha[75][56] = 1'b1; \
	doodle_left_alpha[75][57] = 1'b0; \
	doodle_left_alpha[75][58] = 1'b0; \
	doodle_left_alpha[75][59] = 1'b0; \
	doodle_left_alpha[75][60] = 1'b0; \
	doodle_left_alpha[75][61] = 1'b1; \
	doodle_left_alpha[75][62] = 1'b1; \
	doodle_left_alpha[75][63] = 1'b1; \
	doodle_left_alpha[75][64] = 1'b1; \
	doodle_left_alpha[75][65] = 1'b1; \
	doodle_left_alpha[75][66] = 1'b1; \
	doodle_left_alpha[75][67] = 1'b1; \
	doodle_left_alpha[75][68] = 1'b1; \
	doodle_left_alpha[75][69] = 1'b1; \
	doodle_left_alpha[75][70] = 1'b1; \
	doodle_left_alpha[75][71] = 1'b1; \
	doodle_left_alpha[75][72] = 1'b1; \
	doodle_left_alpha[75][73] = 1'b1; \
	doodle_left_alpha[75][74] = 1'b1; \
	doodle_left_alpha[75][75] = 1'b1; \
	doodle_left_alpha[75][76] = 1'b1; \
	doodle_left_alpha[75][77] = 1'b1; \
	doodle_left_alpha[75][78] = 1'b1; \
	doodle_left_alpha[75][79] = 1'b1; \
	doodle_left_alpha[76][0] = 1'b1; \
	doodle_left_alpha[76][1] = 1'b1; \
	doodle_left_alpha[76][2] = 1'b1; \
	doodle_left_alpha[76][3] = 1'b1; \
	doodle_left_alpha[76][4] = 1'b1; \
	doodle_left_alpha[76][5] = 1'b1; \
	doodle_left_alpha[76][6] = 1'b1; \
	doodle_left_alpha[76][7] = 1'b1; \
	doodle_left_alpha[76][8] = 1'b1; \
	doodle_left_alpha[76][9] = 1'b1; \
	doodle_left_alpha[76][10] = 1'b1; \
	doodle_left_alpha[76][11] = 1'b1; \
	doodle_left_alpha[76][12] = 1'b1; \
	doodle_left_alpha[76][13] = 1'b1; \
	doodle_left_alpha[76][14] = 1'b1; \
	doodle_left_alpha[76][15] = 1'b1; \
	doodle_left_alpha[76][16] = 1'b1; \
	doodle_left_alpha[76][17] = 1'b1; \
	doodle_left_alpha[76][18] = 1'b1; \
	doodle_left_alpha[76][19] = 1'b1; \
	doodle_left_alpha[76][20] = 1'b1; \
	doodle_left_alpha[76][21] = 1'b1; \
	doodle_left_alpha[76][22] = 1'b1; \
	doodle_left_alpha[76][23] = 1'b0; \
	doodle_left_alpha[76][24] = 1'b0; \
	doodle_left_alpha[76][25] = 1'b0; \
	doodle_left_alpha[76][26] = 1'b0; \
	doodle_left_alpha[76][27] = 1'b0; \
	doodle_left_alpha[76][28] = 1'b0; \
	doodle_left_alpha[76][29] = 1'b0; \
	doodle_left_alpha[76][30] = 1'b0; \
	doodle_left_alpha[76][31] = 1'b1; \
	doodle_left_alpha[76][32] = 1'b1; \
	doodle_left_alpha[76][33] = 1'b0; \
	doodle_left_alpha[76][34] = 1'b0; \
	doodle_left_alpha[76][35] = 1'b0; \
	doodle_left_alpha[76][36] = 1'b0; \
	doodle_left_alpha[76][37] = 1'b0; \
	doodle_left_alpha[76][38] = 1'b0; \
	doodle_left_alpha[76][39] = 1'b0; \
	doodle_left_alpha[76][40] = 1'b0; \
	doodle_left_alpha[76][41] = 1'b1; \
	doodle_left_alpha[76][42] = 1'b1; \
	doodle_left_alpha[76][43] = 1'b0; \
	doodle_left_alpha[76][44] = 1'b0; \
	doodle_left_alpha[76][45] = 1'b0; \
	doodle_left_alpha[76][46] = 1'b0; \
	doodle_left_alpha[76][47] = 1'b0; \
	doodle_left_alpha[76][48] = 1'b0; \
	doodle_left_alpha[76][49] = 1'b0; \
	doodle_left_alpha[76][50] = 1'b0; \
	doodle_left_alpha[76][51] = 1'b1; \
	doodle_left_alpha[76][52] = 1'b1; \
	doodle_left_alpha[76][53] = 1'b0; \
	doodle_left_alpha[76][54] = 1'b0; \
	doodle_left_alpha[76][55] = 1'b0; \
	doodle_left_alpha[76][56] = 1'b0; \
	doodle_left_alpha[76][57] = 1'b0; \
	doodle_left_alpha[76][58] = 1'b0; \
	doodle_left_alpha[76][59] = 1'b0; \
	doodle_left_alpha[76][60] = 1'b0; \
	doodle_left_alpha[76][61] = 1'b1; \
	doodle_left_alpha[76][62] = 1'b1; \
	doodle_left_alpha[76][63] = 1'b1; \
	doodle_left_alpha[76][64] = 1'b1; \
	doodle_left_alpha[76][65] = 1'b1; \
	doodle_left_alpha[76][66] = 1'b1; \
	doodle_left_alpha[76][67] = 1'b1; \
	doodle_left_alpha[76][68] = 1'b1; \
	doodle_left_alpha[76][69] = 1'b1; \
	doodle_left_alpha[76][70] = 1'b1; \
	doodle_left_alpha[76][71] = 1'b1; \
	doodle_left_alpha[76][72] = 1'b1; \
	doodle_left_alpha[76][73] = 1'b1; \
	doodle_left_alpha[76][74] = 1'b1; \
	doodle_left_alpha[76][75] = 1'b1; \
	doodle_left_alpha[76][76] = 1'b1; \
	doodle_left_alpha[76][77] = 1'b1; \
	doodle_left_alpha[76][78] = 1'b1; \
	doodle_left_alpha[76][79] = 1'b1; \
	doodle_left_alpha[77][0] = 1'b1; \
	doodle_left_alpha[77][1] = 1'b1; \
	doodle_left_alpha[77][2] = 1'b1; \
	doodle_left_alpha[77][3] = 1'b1; \
	doodle_left_alpha[77][4] = 1'b1; \
	doodle_left_alpha[77][5] = 1'b1; \
	doodle_left_alpha[77][6] = 1'b1; \
	doodle_left_alpha[77][7] = 1'b1; \
	doodle_left_alpha[77][8] = 1'b1; \
	doodle_left_alpha[77][9] = 1'b1; \
	doodle_left_alpha[77][10] = 1'b1; \
	doodle_left_alpha[77][11] = 1'b1; \
	doodle_left_alpha[77][12] = 1'b1; \
	doodle_left_alpha[77][13] = 1'b1; \
	doodle_left_alpha[77][14] = 1'b1; \
	doodle_left_alpha[77][15] = 1'b1; \
	doodle_left_alpha[77][16] = 1'b1; \
	doodle_left_alpha[77][17] = 1'b1; \
	doodle_left_alpha[77][18] = 1'b1; \
	doodle_left_alpha[77][19] = 1'b1; \
	doodle_left_alpha[77][20] = 1'b1; \
	doodle_left_alpha[77][21] = 1'b1; \
	doodle_left_alpha[77][22] = 1'b1; \
	doodle_left_alpha[77][23] = 1'b0; \
	doodle_left_alpha[77][24] = 1'b0; \
	doodle_left_alpha[77][25] = 1'b0; \
	doodle_left_alpha[77][26] = 1'b0; \
	doodle_left_alpha[77][27] = 1'b0; \
	doodle_left_alpha[77][28] = 1'b0; \
	doodle_left_alpha[77][29] = 1'b0; \
	doodle_left_alpha[77][30] = 1'b0; \
	doodle_left_alpha[77][31] = 1'b1; \
	doodle_left_alpha[77][32] = 1'b1; \
	doodle_left_alpha[77][33] = 1'b0; \
	doodle_left_alpha[77][34] = 1'b0; \
	doodle_left_alpha[77][35] = 1'b0; \
	doodle_left_alpha[77][36] = 1'b0; \
	doodle_left_alpha[77][37] = 1'b0; \
	doodle_left_alpha[77][38] = 1'b0; \
	doodle_left_alpha[77][39] = 1'b0; \
	doodle_left_alpha[77][40] = 1'b0; \
	doodle_left_alpha[77][41] = 1'b1; \
	doodle_left_alpha[77][42] = 1'b1; \
	doodle_left_alpha[77][43] = 1'b0; \
	doodle_left_alpha[77][44] = 1'b0; \
	doodle_left_alpha[77][45] = 1'b0; \
	doodle_left_alpha[77][46] = 1'b0; \
	doodle_left_alpha[77][47] = 1'b0; \
	doodle_left_alpha[77][48] = 1'b0; \
	doodle_left_alpha[77][49] = 1'b0; \
	doodle_left_alpha[77][50] = 1'b0; \
	doodle_left_alpha[77][51] = 1'b1; \
	doodle_left_alpha[77][52] = 1'b1; \
	doodle_left_alpha[77][53] = 1'b0; \
	doodle_left_alpha[77][54] = 1'b0; \
	doodle_left_alpha[77][55] = 1'b0; \
	doodle_left_alpha[77][56] = 1'b0; \
	doodle_left_alpha[77][57] = 1'b0; \
	doodle_left_alpha[77][58] = 1'b0; \
	doodle_left_alpha[77][59] = 1'b0; \
	doodle_left_alpha[77][60] = 1'b0; \
	doodle_left_alpha[77][61] = 1'b1; \
	doodle_left_alpha[77][62] = 1'b1; \
	doodle_left_alpha[77][63] = 1'b1; \
	doodle_left_alpha[77][64] = 1'b1; \
	doodle_left_alpha[77][65] = 1'b1; \
	doodle_left_alpha[77][66] = 1'b1; \
	doodle_left_alpha[77][67] = 1'b1; \
	doodle_left_alpha[77][68] = 1'b1; \
	doodle_left_alpha[77][69] = 1'b1; \
	doodle_left_alpha[77][70] = 1'b1; \
	doodle_left_alpha[77][71] = 1'b1; \
	doodle_left_alpha[77][72] = 1'b1; \
	doodle_left_alpha[77][73] = 1'b1; \
	doodle_left_alpha[77][74] = 1'b1; \
	doodle_left_alpha[77][75] = 1'b1; \
	doodle_left_alpha[77][76] = 1'b1; \
	doodle_left_alpha[77][77] = 1'b1; \
	doodle_left_alpha[77][78] = 1'b1; \
	doodle_left_alpha[77][79] = 1'b1; \
	doodle_left_alpha[78][0] = 1'b1; \
	doodle_left_alpha[78][1] = 1'b1; \
	doodle_left_alpha[78][2] = 1'b1; \
	doodle_left_alpha[78][3] = 1'b1; \
	doodle_left_alpha[78][4] = 1'b1; \
	doodle_left_alpha[78][5] = 1'b1; \
	doodle_left_alpha[78][6] = 1'b1; \
	doodle_left_alpha[78][7] = 1'b1; \
	doodle_left_alpha[78][8] = 1'b1; \
	doodle_left_alpha[78][9] = 1'b1; \
	doodle_left_alpha[78][10] = 1'b1; \
	doodle_left_alpha[78][11] = 1'b1; \
	doodle_left_alpha[78][12] = 1'b1; \
	doodle_left_alpha[78][13] = 1'b1; \
	doodle_left_alpha[78][14] = 1'b1; \
	doodle_left_alpha[78][15] = 1'b1; \
	doodle_left_alpha[78][16] = 1'b1; \
	doodle_left_alpha[78][17] = 1'b1; \
	doodle_left_alpha[78][18] = 1'b1; \
	doodle_left_alpha[78][19] = 1'b1; \
	doodle_left_alpha[78][20] = 1'b1; \
	doodle_left_alpha[78][21] = 1'b1; \
	doodle_left_alpha[78][22] = 1'b1; \
	doodle_left_alpha[78][23] = 1'b0; \
	doodle_left_alpha[78][24] = 1'b0; \
	doodle_left_alpha[78][25] = 1'b0; \
	doodle_left_alpha[78][26] = 1'b0; \
	doodle_left_alpha[78][27] = 1'b0; \
	doodle_left_alpha[78][28] = 1'b0; \
	doodle_left_alpha[78][29] = 1'b0; \
	doodle_left_alpha[78][30] = 1'b0; \
	doodle_left_alpha[78][31] = 1'b1; \
	doodle_left_alpha[78][32] = 1'b1; \
	doodle_left_alpha[78][33] = 1'b0; \
	doodle_left_alpha[78][34] = 1'b0; \
	doodle_left_alpha[78][35] = 1'b0; \
	doodle_left_alpha[78][36] = 1'b0; \
	doodle_left_alpha[78][37] = 1'b0; \
	doodle_left_alpha[78][38] = 1'b0; \
	doodle_left_alpha[78][39] = 1'b0; \
	doodle_left_alpha[78][40] = 1'b0; \
	doodle_left_alpha[78][41] = 1'b1; \
	doodle_left_alpha[78][42] = 1'b1; \
	doodle_left_alpha[78][43] = 1'b0; \
	doodle_left_alpha[78][44] = 1'b0; \
	doodle_left_alpha[78][45] = 1'b0; \
	doodle_left_alpha[78][46] = 1'b0; \
	doodle_left_alpha[78][47] = 1'b0; \
	doodle_left_alpha[78][48] = 1'b0; \
	doodle_left_alpha[78][49] = 1'b0; \
	doodle_left_alpha[78][50] = 1'b0; \
	doodle_left_alpha[78][51] = 1'b1; \
	doodle_left_alpha[78][52] = 1'b1; \
	doodle_left_alpha[78][53] = 1'b0; \
	doodle_left_alpha[78][54] = 1'b0; \
	doodle_left_alpha[78][55] = 1'b0; \
	doodle_left_alpha[78][56] = 1'b0; \
	doodle_left_alpha[78][57] = 1'b0; \
	doodle_left_alpha[78][58] = 1'b0; \
	doodle_left_alpha[78][59] = 1'b0; \
	doodle_left_alpha[78][60] = 1'b0; \
	doodle_left_alpha[78][61] = 1'b1; \
	doodle_left_alpha[78][62] = 1'b1; \
	doodle_left_alpha[78][63] = 1'b1; \
	doodle_left_alpha[78][64] = 1'b1; \
	doodle_left_alpha[78][65] = 1'b1; \
	doodle_left_alpha[78][66] = 1'b1; \
	doodle_left_alpha[78][67] = 1'b1; \
	doodle_left_alpha[78][68] = 1'b1; \
	doodle_left_alpha[78][69] = 1'b1; \
	doodle_left_alpha[78][70] = 1'b1; \
	doodle_left_alpha[78][71] = 1'b1; \
	doodle_left_alpha[78][72] = 1'b1; \
	doodle_left_alpha[78][73] = 1'b1; \
	doodle_left_alpha[78][74] = 1'b1; \
	doodle_left_alpha[78][75] = 1'b1; \
	doodle_left_alpha[78][76] = 1'b1; \
	doodle_left_alpha[78][77] = 1'b1; \
	doodle_left_alpha[78][78] = 1'b1; \
	doodle_left_alpha[78][79] = 1'b1; \
	doodle_left_alpha[79][0] = 1'b1; \
	doodle_left_alpha[79][1] = 1'b1; \
	doodle_left_alpha[79][2] = 1'b1; \
	doodle_left_alpha[79][3] = 1'b1; \
	doodle_left_alpha[79][4] = 1'b1; \
	doodle_left_alpha[79][5] = 1'b1; \
	doodle_left_alpha[79][6] = 1'b1; \
	doodle_left_alpha[79][7] = 1'b1; \
	doodle_left_alpha[79][8] = 1'b1; \
	doodle_left_alpha[79][9] = 1'b1; \
	doodle_left_alpha[79][10] = 1'b1; \
	doodle_left_alpha[79][11] = 1'b1; \
	doodle_left_alpha[79][12] = 1'b1; \
	doodle_left_alpha[79][13] = 1'b1; \
	doodle_left_alpha[79][14] = 1'b1; \
	doodle_left_alpha[79][15] = 1'b1; \
	doodle_left_alpha[79][16] = 1'b1; \
	doodle_left_alpha[79][17] = 1'b1; \
	doodle_left_alpha[79][18] = 1'b1; \
	doodle_left_alpha[79][19] = 1'b1; \
	doodle_left_alpha[79][20] = 1'b1; \
	doodle_left_alpha[79][21] = 1'b1; \
	doodle_left_alpha[79][22] = 1'b1; \
	doodle_left_alpha[79][23] = 1'b0; \
	doodle_left_alpha[79][24] = 1'b0; \
	doodle_left_alpha[79][25] = 1'b0; \
	doodle_left_alpha[79][26] = 1'b0; \
	doodle_left_alpha[79][27] = 1'b0; \
	doodle_left_alpha[79][28] = 1'b0; \
	doodle_left_alpha[79][29] = 1'b0; \
	doodle_left_alpha[79][30] = 1'b0; \
	doodle_left_alpha[79][31] = 1'b1; \
	doodle_left_alpha[79][32] = 1'b1; \
	doodle_left_alpha[79][33] = 1'b0; \
	doodle_left_alpha[79][34] = 1'b0; \
	doodle_left_alpha[79][35] = 1'b0; \
	doodle_left_alpha[79][36] = 1'b0; \
	doodle_left_alpha[79][37] = 1'b0; \
	doodle_left_alpha[79][38] = 1'b0; \
	doodle_left_alpha[79][39] = 1'b0; \
	doodle_left_alpha[79][40] = 1'b0; \
	doodle_left_alpha[79][41] = 1'b1; \
	doodle_left_alpha[79][42] = 1'b1; \
	doodle_left_alpha[79][43] = 1'b0; \
	doodle_left_alpha[79][44] = 1'b0; \
	doodle_left_alpha[79][45] = 1'b0; \
	doodle_left_alpha[79][46] = 1'b0; \
	doodle_left_alpha[79][47] = 1'b0; \
	doodle_left_alpha[79][48] = 1'b0; \
	doodle_left_alpha[79][49] = 1'b0; \
	doodle_left_alpha[79][50] = 1'b0; \
	doodle_left_alpha[79][51] = 1'b1; \
	doodle_left_alpha[79][52] = 1'b1; \
	doodle_left_alpha[79][53] = 1'b0; \
	doodle_left_alpha[79][54] = 1'b0; \
	doodle_left_alpha[79][55] = 1'b0; \
	doodle_left_alpha[79][56] = 1'b0; \
	doodle_left_alpha[79][57] = 1'b0; \
	doodle_left_alpha[79][58] = 1'b0; \
	doodle_left_alpha[79][59] = 1'b0; \
	doodle_left_alpha[79][60] = 1'b0; \
	doodle_left_alpha[79][61] = 1'b1; \
	doodle_left_alpha[79][62] = 1'b1; \
	doodle_left_alpha[79][63] = 1'b1; \
	doodle_left_alpha[79][64] = 1'b1; \
	doodle_left_alpha[79][65] = 1'b1; \
	doodle_left_alpha[79][66] = 1'b1; \
	doodle_left_alpha[79][67] = 1'b1; \
	doodle_left_alpha[79][68] = 1'b1; \
	doodle_left_alpha[79][69] = 1'b1; \
	doodle_left_alpha[79][70] = 1'b1; \
	doodle_left_alpha[79][71] = 1'b1; \
	doodle_left_alpha[79][72] = 1'b1; \
	doodle_left_alpha[79][73] = 1'b1; \
	doodle_left_alpha[79][74] = 1'b1; \
	doodle_left_alpha[79][75] = 1'b1; \
	doodle_left_alpha[79][76] = 1'b1; \
	doodle_left_alpha[79][77] = 1'b1; \
	doodle_left_alpha[79][78] = 1'b1; \
	doodle_left_alpha[79][79] = 1'b1; \
end

`endif // INITIAL_DOODLE_LEFT
