module platforms(
	input clk,
	input rst,
	
	output logic [9:0] led,

	input [10:0] beam_x,
	input [9:0] beam_y,

	output logic signed [92:0][1:0][10:0] platforms,
	output logic [92:0] platform_activation,
	
	output logic [2:0][3:0] color,
	output logic is_transparent
);

logic [29:0][99:0][2:0][3:0] green_platform_texture;
logic [29:0][99:0] green_platform_transparency_texture;
logic [92:0] draw;
logic [6:0] here_platform_was_generated;

/*assign platforms[0][1] = 342;
assign platforms[0][0] = -10;
assign led[0] = platforms[0][0] < 0;*/

logic [15:0] random_sides;
random_sonya_coin sonya_coin(
	.clk(clk),
	.rst(rst),
	
	.fibonacci_LSFR(random_sides)
);

//localparam [92:0] random_start = 93'b000000000000000000000000000000000010000100000001010000000010000000001000000000000110000100001;
localparam [92:0] random_start = 93'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
always_ff @ (posedge clk) begin
	if (rst) begin
		for (int i = 0; i < 31; i++)
			for (int j = 0; j < 3; j++) begin
				platforms[i * 3 + j][0] <= -162 + i * 30;
				platforms[i * 3 + j][1] <= 342 + j * 114;	
			end
		// random activation (6 fors + control)
		for (int j = 0; j < 7; j++)
			for (int i = 0; i < (j < 6 ? 15 : 3); i++) begin
				if (j * 15 + i > 74) platform_activation[j * 15 + i] <= 0;
				else if (i == (j < 6 ? 14 : 2) && ~here_platform_was_generated[j])
					platform_activation[j * 15 + i] <= 0;
				else begin
					platform_activation[j * 15 + i] <= random_start[j * 15 + i];
					if (i == 0) here_platform_was_generated[j] <= platform_activation[j * 15 + i];
					else here_platform_was_generated[j] <= here_platform_was_generated[j] || platform_activation[j * 15 + i];
				end
			end
	end else begin
		
	end
end

genvar i;
generate 
	for (i = 0; i < 93; i++) begin: name
		assign draw[i] =  $signed(platforms[i][1]) <= $signed(beam_x) && $signed(beam_x) <= $signed(platforms[i][1]) + 100 - 1
			&& $signed(platforms[i][0]) <= $signed(11'(beam_y)) && $signed(11'(beam_y)) <= $signed(platforms[i][0]) + 30 - 1 && platform_activation[i];
	end
endgenerate

always_ff @(posedge clk) begin
	for (int i = 0; i < 93; i++) begin 
		if (draw[i]) begin 
			color[0] = green_platform_texture[beam_y - platforms[i][0]][beam_x - platforms[i][1]][0];
			color[1] = green_platform_texture[beam_y - platforms[i][0]][beam_x - platforms[i][1]][1];
			color[2] = green_platform_texture[beam_y - platforms[i][0]][beam_x - platforms[i][1]][2];
			is_transparent = green_platform_transparency_texture[beam_y - platforms[i][0]][beam_x - platforms[i][1]];
		end 
	end
	if (~|draw) begin 
		is_transparent = 1; 
		color = '1;
	end
end

always_comb begin
	green_platform_texture[0][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[0][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[1][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[2][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[3][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[4][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[5][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[6][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[7][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[8][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[9][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[10][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[10][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[11][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[11][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[12][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[12][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[13][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[13][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[14][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[14][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[15][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[15][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[16][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[16][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[17][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[17][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[18][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[18][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][10] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][11] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][12] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][13] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][14] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][15] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][16] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][17] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][18] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][19] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][20] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][21] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][22] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][23] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][24] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][25] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][26] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][27] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][28] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][29] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][30] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][31] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][32] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][33] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][34] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][35] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][36] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][37] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][38] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][39] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][40] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][41] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][42] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][43] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][44] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][45] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][46] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][47] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][48] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][49] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][50] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][51] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][52] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][53] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][54] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][55] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][56] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][57] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][58] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][59] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][60] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][61] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][62] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][63] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][64] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][65] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][66] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][67] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][68] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][69] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][70] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][71] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][72] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][73] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][74] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][75] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][76] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][77] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][78] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][79] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][80] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][81] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][82] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][83] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][84] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][85] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][86] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][87] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][88] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][89] = {4'b0, 4'b1111, 4'b0};	green_platform_texture[19][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[19][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[20][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[21][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[22][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[23][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[24][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[25][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[26][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[27][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[28][99] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][0] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][1] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][2] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][3] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][4] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][5] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][6] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][7] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][8] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][9] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][10] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][11] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][12] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][13] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][14] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][15] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][16] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][17] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][18] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][19] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][20] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][21] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][22] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][23] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][24] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][25] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][26] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][27] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][28] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][29] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][30] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][31] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][32] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][33] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][34] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][35] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][36] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][37] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][38] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][39] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][40] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][41] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][42] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][43] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][44] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][45] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][46] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][47] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][48] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][49] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][50] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][51] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][52] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][53] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][54] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][55] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][56] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][57] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][58] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][59] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][60] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][61] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][62] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][63] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][64] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][65] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][66] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][67] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][68] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][69] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][70] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][71] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][72] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][73] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][74] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][75] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][76] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][77] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][78] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][79] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][80] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][81] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][82] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][83] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][84] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][85] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][86] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][87] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][88] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][89] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][90] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][91] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][92] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][93] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][94] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][95] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][96] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][97] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][98] = {4'b0, 4'b0, 4'b0};	green_platform_texture[29][99] = {4'b0, 4'b0, 4'b0};
	green_platform_transparency_texture[0][0] = 1;	green_platform_transparency_texture[0][1] = 1;	green_platform_transparency_texture[0][2] = 1;	green_platform_transparency_texture[0][3] = 1;	green_platform_transparency_texture[0][4] = 1;	green_platform_transparency_texture[0][5] = 1;	green_platform_transparency_texture[0][6] = 1;	green_platform_transparency_texture[0][7] = 1;	green_platform_transparency_texture[0][8] = 1;	green_platform_transparency_texture[0][9] = 1;	green_platform_transparency_texture[0][10] = 1;	green_platform_transparency_texture[0][11] = 1;	green_platform_transparency_texture[0][12] = 1;	green_platform_transparency_texture[0][13] = 1;	green_platform_transparency_texture[0][14] = 1;	green_platform_transparency_texture[0][15] = 1;	green_platform_transparency_texture[0][16] = 1;	green_platform_transparency_texture[0][17] = 1;	green_platform_transparency_texture[0][18] = 1;	green_platform_transparency_texture[0][19] = 1;	green_platform_transparency_texture[0][20] = 1;	green_platform_transparency_texture[0][21] = 1;	green_platform_transparency_texture[0][22] = 1;	green_platform_transparency_texture[0][23] = 1;	green_platform_transparency_texture[0][24] = 1;	green_platform_transparency_texture[0][25] = 1;	green_platform_transparency_texture[0][26] = 1;	green_platform_transparency_texture[0][27] = 1;	green_platform_transparency_texture[0][28] = 1;	green_platform_transparency_texture[0][29] = 1;	green_platform_transparency_texture[0][30] = 1;	green_platform_transparency_texture[0][31] = 1;	green_platform_transparency_texture[0][32] = 1;	green_platform_transparency_texture[0][33] = 1;	green_platform_transparency_texture[0][34] = 1;	green_platform_transparency_texture[0][35] = 1;	green_platform_transparency_texture[0][36] = 1;	green_platform_transparency_texture[0][37] = 1;	green_platform_transparency_texture[0][38] = 1;	green_platform_transparency_texture[0][39] = 1;	green_platform_transparency_texture[0][40] = 1;	green_platform_transparency_texture[0][41] = 1;	green_platform_transparency_texture[0][42] = 1;	green_platform_transparency_texture[0][43] = 1;	green_platform_transparency_texture[0][44] = 1;	green_platform_transparency_texture[0][45] = 1;	green_platform_transparency_texture[0][46] = 1;	green_platform_transparency_texture[0][47] = 1;	green_platform_transparency_texture[0][48] = 1;	green_platform_transparency_texture[0][49] = 1;	green_platform_transparency_texture[0][50] = 1;	green_platform_transparency_texture[0][51] = 1;	green_platform_transparency_texture[0][52] = 1;	green_platform_transparency_texture[0][53] = 1;	green_platform_transparency_texture[0][54] = 1;	green_platform_transparency_texture[0][55] = 1;	green_platform_transparency_texture[0][56] = 1;	green_platform_transparency_texture[0][57] = 1;	green_platform_transparency_texture[0][58] = 1;	green_platform_transparency_texture[0][59] = 1;	green_platform_transparency_texture[0][60] = 1;	green_platform_transparency_texture[0][61] = 1;	green_platform_transparency_texture[0][62] = 1;	green_platform_transparency_texture[0][63] = 1;	green_platform_transparency_texture[0][64] = 1;	green_platform_transparency_texture[0][65] = 1;	green_platform_transparency_texture[0][66] = 1;	green_platform_transparency_texture[0][67] = 1;	green_platform_transparency_texture[0][68] = 1;	green_platform_transparency_texture[0][69] = 1;	green_platform_transparency_texture[0][70] = 1;	green_platform_transparency_texture[0][71] = 1;	green_platform_transparency_texture[0][72] = 1;	green_platform_transparency_texture[0][73] = 1;	green_platform_transparency_texture[0][74] = 1;	green_platform_transparency_texture[0][75] = 1;	green_platform_transparency_texture[0][76] = 1;	green_platform_transparency_texture[0][77] = 1;	green_platform_transparency_texture[0][78] = 1;	green_platform_transparency_texture[0][79] = 1;	green_platform_transparency_texture[0][80] = 1;	green_platform_transparency_texture[0][81] = 1;	green_platform_transparency_texture[0][82] = 1;	green_platform_transparency_texture[0][83] = 1;	green_platform_transparency_texture[0][84] = 1;	green_platform_transparency_texture[0][85] = 1;	green_platform_transparency_texture[0][86] = 1;	green_platform_transparency_texture[0][87] = 1;	green_platform_transparency_texture[0][88] = 1;	green_platform_transparency_texture[0][89] = 1;	green_platform_transparency_texture[0][90] = 1;	green_platform_transparency_texture[0][91] = 1;	green_platform_transparency_texture[0][92] = 1;	green_platform_transparency_texture[0][93] = 1;	green_platform_transparency_texture[0][94] = 1;	green_platform_transparency_texture[0][95] = 1;	green_platform_transparency_texture[0][96] = 1;	green_platform_transparency_texture[0][97] = 1;	green_platform_transparency_texture[0][98] = 1;	green_platform_transparency_texture[0][99] = 1;	green_platform_transparency_texture[1][0] = 1;	green_platform_transparency_texture[1][1] = 1;	green_platform_transparency_texture[1][2] = 1;	green_platform_transparency_texture[1][3] = 1;	green_platform_transparency_texture[1][4] = 1;	green_platform_transparency_texture[1][5] = 1;	green_platform_transparency_texture[1][6] = 1;	green_platform_transparency_texture[1][7] = 1;	green_platform_transparency_texture[1][8] = 1;	green_platform_transparency_texture[1][9] = 1;	green_platform_transparency_texture[1][10] = 1;	green_platform_transparency_texture[1][11] = 1;	green_platform_transparency_texture[1][12] = 1;	green_platform_transparency_texture[1][13] = 1;	green_platform_transparency_texture[1][14] = 1;	green_platform_transparency_texture[1][15] = 1;	green_platform_transparency_texture[1][16] = 1;	green_platform_transparency_texture[1][17] = 1;	green_platform_transparency_texture[1][18] = 1;	green_platform_transparency_texture[1][19] = 1;	green_platform_transparency_texture[1][20] = 1;	green_platform_transparency_texture[1][21] = 1;	green_platform_transparency_texture[1][22] = 1;	green_platform_transparency_texture[1][23] = 1;	green_platform_transparency_texture[1][24] = 1;	green_platform_transparency_texture[1][25] = 1;	green_platform_transparency_texture[1][26] = 1;	green_platform_transparency_texture[1][27] = 1;	green_platform_transparency_texture[1][28] = 1;	green_platform_transparency_texture[1][29] = 1;	green_platform_transparency_texture[1][30] = 1;	green_platform_transparency_texture[1][31] = 1;	green_platform_transparency_texture[1][32] = 1;	green_platform_transparency_texture[1][33] = 1;	green_platform_transparency_texture[1][34] = 1;	green_platform_transparency_texture[1][35] = 1;	green_platform_transparency_texture[1][36] = 1;	green_platform_transparency_texture[1][37] = 1;	green_platform_transparency_texture[1][38] = 1;	green_platform_transparency_texture[1][39] = 1;	green_platform_transparency_texture[1][40] = 1;	green_platform_transparency_texture[1][41] = 1;	green_platform_transparency_texture[1][42] = 1;	green_platform_transparency_texture[1][43] = 1;	green_platform_transparency_texture[1][44] = 1;	green_platform_transparency_texture[1][45] = 1;	green_platform_transparency_texture[1][46] = 1;	green_platform_transparency_texture[1][47] = 1;	green_platform_transparency_texture[1][48] = 1;	green_platform_transparency_texture[1][49] = 1;	green_platform_transparency_texture[1][50] = 1;	green_platform_transparency_texture[1][51] = 1;	green_platform_transparency_texture[1][52] = 1;	green_platform_transparency_texture[1][53] = 1;	green_platform_transparency_texture[1][54] = 1;	green_platform_transparency_texture[1][55] = 1;	green_platform_transparency_texture[1][56] = 1;	green_platform_transparency_texture[1][57] = 1;	green_platform_transparency_texture[1][58] = 1;	green_platform_transparency_texture[1][59] = 1;	green_platform_transparency_texture[1][60] = 1;	green_platform_transparency_texture[1][61] = 1;	green_platform_transparency_texture[1][62] = 1;	green_platform_transparency_texture[1][63] = 1;	green_platform_transparency_texture[1][64] = 1;	green_platform_transparency_texture[1][65] = 1;	green_platform_transparency_texture[1][66] = 1;	green_platform_transparency_texture[1][67] = 1;	green_platform_transparency_texture[1][68] = 1;	green_platform_transparency_texture[1][69] = 1;	green_platform_transparency_texture[1][70] = 1;	green_platform_transparency_texture[1][71] = 1;	green_platform_transparency_texture[1][72] = 1;	green_platform_transparency_texture[1][73] = 1;	green_platform_transparency_texture[1][74] = 1;	green_platform_transparency_texture[1][75] = 1;	green_platform_transparency_texture[1][76] = 1;	green_platform_transparency_texture[1][77] = 1;	green_platform_transparency_texture[1][78] = 1;	green_platform_transparency_texture[1][79] = 1;	green_platform_transparency_texture[1][80] = 1;	green_platform_transparency_texture[1][81] = 1;	green_platform_transparency_texture[1][82] = 1;	green_platform_transparency_texture[1][83] = 1;	green_platform_transparency_texture[1][84] = 1;	green_platform_transparency_texture[1][85] = 1;	green_platform_transparency_texture[1][86] = 1;	green_platform_transparency_texture[1][87] = 1;	green_platform_transparency_texture[1][88] = 1;	green_platform_transparency_texture[1][89] = 1;	green_platform_transparency_texture[1][90] = 1;	green_platform_transparency_texture[1][91] = 1;	green_platform_transparency_texture[1][92] = 1;	green_platform_transparency_texture[1][93] = 1;	green_platform_transparency_texture[1][94] = 1;	green_platform_transparency_texture[1][95] = 1;	green_platform_transparency_texture[1][96] = 1;	green_platform_transparency_texture[1][97] = 1;	green_platform_transparency_texture[1][98] = 1;	green_platform_transparency_texture[1][99] = 1;	green_platform_transparency_texture[2][0] = 1;	green_platform_transparency_texture[2][1] = 1;	green_platform_transparency_texture[2][2] = 1;	green_platform_transparency_texture[2][3] = 1;	green_platform_transparency_texture[2][4] = 1;	green_platform_transparency_texture[2][5] = 1;	green_platform_transparency_texture[2][6] = 1;	green_platform_transparency_texture[2][7] = 1;	green_platform_transparency_texture[2][8] = 1;	green_platform_transparency_texture[2][9] = 1;	green_platform_transparency_texture[2][10] = 1;	green_platform_transparency_texture[2][11] = 1;	green_platform_transparency_texture[2][12] = 1;	green_platform_transparency_texture[2][13] = 1;	green_platform_transparency_texture[2][14] = 1;	green_platform_transparency_texture[2][15] = 1;	green_platform_transparency_texture[2][16] = 1;	green_platform_transparency_texture[2][17] = 1;	green_platform_transparency_texture[2][18] = 1;	green_platform_transparency_texture[2][19] = 1;	green_platform_transparency_texture[2][20] = 1;	green_platform_transparency_texture[2][21] = 1;	green_platform_transparency_texture[2][22] = 1;	green_platform_transparency_texture[2][23] = 1;	green_platform_transparency_texture[2][24] = 1;	green_platform_transparency_texture[2][25] = 1;	green_platform_transparency_texture[2][26] = 1;	green_platform_transparency_texture[2][27] = 1;	green_platform_transparency_texture[2][28] = 1;	green_platform_transparency_texture[2][29] = 1;	green_platform_transparency_texture[2][30] = 1;	green_platform_transparency_texture[2][31] = 1;	green_platform_transparency_texture[2][32] = 1;	green_platform_transparency_texture[2][33] = 1;	green_platform_transparency_texture[2][34] = 1;	green_platform_transparency_texture[2][35] = 1;	green_platform_transparency_texture[2][36] = 1;	green_platform_transparency_texture[2][37] = 1;	green_platform_transparency_texture[2][38] = 1;	green_platform_transparency_texture[2][39] = 1;	green_platform_transparency_texture[2][40] = 1;	green_platform_transparency_texture[2][41] = 1;	green_platform_transparency_texture[2][42] = 1;	green_platform_transparency_texture[2][43] = 1;	green_platform_transparency_texture[2][44] = 1;	green_platform_transparency_texture[2][45] = 1;	green_platform_transparency_texture[2][46] = 1;	green_platform_transparency_texture[2][47] = 1;	green_platform_transparency_texture[2][48] = 1;	green_platform_transparency_texture[2][49] = 1;	green_platform_transparency_texture[2][50] = 1;	green_platform_transparency_texture[2][51] = 1;	green_platform_transparency_texture[2][52] = 1;	green_platform_transparency_texture[2][53] = 1;	green_platform_transparency_texture[2][54] = 1;	green_platform_transparency_texture[2][55] = 1;	green_platform_transparency_texture[2][56] = 1;	green_platform_transparency_texture[2][57] = 1;	green_platform_transparency_texture[2][58] = 1;	green_platform_transparency_texture[2][59] = 1;	green_platform_transparency_texture[2][60] = 1;	green_platform_transparency_texture[2][61] = 1;	green_platform_transparency_texture[2][62] = 1;	green_platform_transparency_texture[2][63] = 1;	green_platform_transparency_texture[2][64] = 1;	green_platform_transparency_texture[2][65] = 1;	green_platform_transparency_texture[2][66] = 1;	green_platform_transparency_texture[2][67] = 1;	green_platform_transparency_texture[2][68] = 1;	green_platform_transparency_texture[2][69] = 1;	green_platform_transparency_texture[2][70] = 1;	green_platform_transparency_texture[2][71] = 1;	green_platform_transparency_texture[2][72] = 1;	green_platform_transparency_texture[2][73] = 1;	green_platform_transparency_texture[2][74] = 1;	green_platform_transparency_texture[2][75] = 1;	green_platform_transparency_texture[2][76] = 1;	green_platform_transparency_texture[2][77] = 1;	green_platform_transparency_texture[2][78] = 1;	green_platform_transparency_texture[2][79] = 1;	green_platform_transparency_texture[2][80] = 1;	green_platform_transparency_texture[2][81] = 1;	green_platform_transparency_texture[2][82] = 1;	green_platform_transparency_texture[2][83] = 1;	green_platform_transparency_texture[2][84] = 1;	green_platform_transparency_texture[2][85] = 1;	green_platform_transparency_texture[2][86] = 1;	green_platform_transparency_texture[2][87] = 1;	green_platform_transparency_texture[2][88] = 1;	green_platform_transparency_texture[2][89] = 1;	green_platform_transparency_texture[2][90] = 1;	green_platform_transparency_texture[2][91] = 1;	green_platform_transparency_texture[2][92] = 1;	green_platform_transparency_texture[2][93] = 1;	green_platform_transparency_texture[2][94] = 1;	green_platform_transparency_texture[2][95] = 1;	green_platform_transparency_texture[2][96] = 1;	green_platform_transparency_texture[2][97] = 1;	green_platform_transparency_texture[2][98] = 1;	green_platform_transparency_texture[2][99] = 1;	green_platform_transparency_texture[3][0] = 1;	green_platform_transparency_texture[3][1] = 1;	green_platform_transparency_texture[3][2] = 1;	green_platform_transparency_texture[3][3] = 1;	green_platform_transparency_texture[3][4] = 1;	green_platform_transparency_texture[3][5] = 1;	green_platform_transparency_texture[3][6] = 1;	green_platform_transparency_texture[3][7] = 1;	green_platform_transparency_texture[3][8] = 1;	green_platform_transparency_texture[3][9] = 1;	green_platform_transparency_texture[3][10] = 1;	green_platform_transparency_texture[3][11] = 1;	green_platform_transparency_texture[3][12] = 1;	green_platform_transparency_texture[3][13] = 1;	green_platform_transparency_texture[3][14] = 1;	green_platform_transparency_texture[3][15] = 1;	green_platform_transparency_texture[3][16] = 1;	green_platform_transparency_texture[3][17] = 1;	green_platform_transparency_texture[3][18] = 1;	green_platform_transparency_texture[3][19] = 1;	green_platform_transparency_texture[3][20] = 1;	green_platform_transparency_texture[3][21] = 1;	green_platform_transparency_texture[3][22] = 1;	green_platform_transparency_texture[3][23] = 1;	green_platform_transparency_texture[3][24] = 1;	green_platform_transparency_texture[3][25] = 1;	green_platform_transparency_texture[3][26] = 1;	green_platform_transparency_texture[3][27] = 1;	green_platform_transparency_texture[3][28] = 1;	green_platform_transparency_texture[3][29] = 1;	green_platform_transparency_texture[3][30] = 1;	green_platform_transparency_texture[3][31] = 1;	green_platform_transparency_texture[3][32] = 1;	green_platform_transparency_texture[3][33] = 1;	green_platform_transparency_texture[3][34] = 1;	green_platform_transparency_texture[3][35] = 1;	green_platform_transparency_texture[3][36] = 1;	green_platform_transparency_texture[3][37] = 1;	green_platform_transparency_texture[3][38] = 1;	green_platform_transparency_texture[3][39] = 1;	green_platform_transparency_texture[3][40] = 1;	green_platform_transparency_texture[3][41] = 1;	green_platform_transparency_texture[3][42] = 1;	green_platform_transparency_texture[3][43] = 1;	green_platform_transparency_texture[3][44] = 1;	green_platform_transparency_texture[3][45] = 1;	green_platform_transparency_texture[3][46] = 1;	green_platform_transparency_texture[3][47] = 1;	green_platform_transparency_texture[3][48] = 1;	green_platform_transparency_texture[3][49] = 1;	green_platform_transparency_texture[3][50] = 1;	green_platform_transparency_texture[3][51] = 1;	green_platform_transparency_texture[3][52] = 1;	green_platform_transparency_texture[3][53] = 1;	green_platform_transparency_texture[3][54] = 1;	green_platform_transparency_texture[3][55] = 1;	green_platform_transparency_texture[3][56] = 1;	green_platform_transparency_texture[3][57] = 1;	green_platform_transparency_texture[3][58] = 1;	green_platform_transparency_texture[3][59] = 1;	green_platform_transparency_texture[3][60] = 1;	green_platform_transparency_texture[3][61] = 1;	green_platform_transparency_texture[3][62] = 1;	green_platform_transparency_texture[3][63] = 1;	green_platform_transparency_texture[3][64] = 1;	green_platform_transparency_texture[3][65] = 1;	green_platform_transparency_texture[3][66] = 1;	green_platform_transparency_texture[3][67] = 1;	green_platform_transparency_texture[3][68] = 1;	green_platform_transparency_texture[3][69] = 1;	green_platform_transparency_texture[3][70] = 1;	green_platform_transparency_texture[3][71] = 1;	green_platform_transparency_texture[3][72] = 1;	green_platform_transparency_texture[3][73] = 1;	green_platform_transparency_texture[3][74] = 1;	green_platform_transparency_texture[3][75] = 1;	green_platform_transparency_texture[3][76] = 1;	green_platform_transparency_texture[3][77] = 1;	green_platform_transparency_texture[3][78] = 1;	green_platform_transparency_texture[3][79] = 1;	green_platform_transparency_texture[3][80] = 1;	green_platform_transparency_texture[3][81] = 1;	green_platform_transparency_texture[3][82] = 1;	green_platform_transparency_texture[3][83] = 1;	green_platform_transparency_texture[3][84] = 1;	green_platform_transparency_texture[3][85] = 1;	green_platform_transparency_texture[3][86] = 1;	green_platform_transparency_texture[3][87] = 1;	green_platform_transparency_texture[3][88] = 1;	green_platform_transparency_texture[3][89] = 1;	green_platform_transparency_texture[3][90] = 1;	green_platform_transparency_texture[3][91] = 1;	green_platform_transparency_texture[3][92] = 1;	green_platform_transparency_texture[3][93] = 1;	green_platform_transparency_texture[3][94] = 1;	green_platform_transparency_texture[3][95] = 1;	green_platform_transparency_texture[3][96] = 1;	green_platform_transparency_texture[3][97] = 1;	green_platform_transparency_texture[3][98] = 1;	green_platform_transparency_texture[3][99] = 1;	green_platform_transparency_texture[4][0] = 1;	green_platform_transparency_texture[4][1] = 1;	green_platform_transparency_texture[4][2] = 1;	green_platform_transparency_texture[4][3] = 1;	green_platform_transparency_texture[4][4] = 1;	green_platform_transparency_texture[4][5] = 1;	green_platform_transparency_texture[4][6] = 1;	green_platform_transparency_texture[4][7] = 1;	green_platform_transparency_texture[4][8] = 1;	green_platform_transparency_texture[4][9] = 1;	green_platform_transparency_texture[4][10] = 1;	green_platform_transparency_texture[4][11] = 1;	green_platform_transparency_texture[4][12] = 1;	green_platform_transparency_texture[4][13] = 1;	green_platform_transparency_texture[4][14] = 1;	green_platform_transparency_texture[4][15] = 1;	green_platform_transparency_texture[4][16] = 1;	green_platform_transparency_texture[4][17] = 1;	green_platform_transparency_texture[4][18] = 1;	green_platform_transparency_texture[4][19] = 1;	green_platform_transparency_texture[4][20] = 1;	green_platform_transparency_texture[4][21] = 1;	green_platform_transparency_texture[4][22] = 1;	green_platform_transparency_texture[4][23] = 1;	green_platform_transparency_texture[4][24] = 1;	green_platform_transparency_texture[4][25] = 1;	green_platform_transparency_texture[4][26] = 1;	green_platform_transparency_texture[4][27] = 1;	green_platform_transparency_texture[4][28] = 1;	green_platform_transparency_texture[4][29] = 1;	green_platform_transparency_texture[4][30] = 1;	green_platform_transparency_texture[4][31] = 1;	green_platform_transparency_texture[4][32] = 1;	green_platform_transparency_texture[4][33] = 1;	green_platform_transparency_texture[4][34] = 1;	green_platform_transparency_texture[4][35] = 1;	green_platform_transparency_texture[4][36] = 1;	green_platform_transparency_texture[4][37] = 1;	green_platform_transparency_texture[4][38] = 1;	green_platform_transparency_texture[4][39] = 1;	green_platform_transparency_texture[4][40] = 1;	green_platform_transparency_texture[4][41] = 1;	green_platform_transparency_texture[4][42] = 1;	green_platform_transparency_texture[4][43] = 1;	green_platform_transparency_texture[4][44] = 1;	green_platform_transparency_texture[4][45] = 1;	green_platform_transparency_texture[4][46] = 1;	green_platform_transparency_texture[4][47] = 1;	green_platform_transparency_texture[4][48] = 1;	green_platform_transparency_texture[4][49] = 1;	green_platform_transparency_texture[4][50] = 1;	green_platform_transparency_texture[4][51] = 1;	green_platform_transparency_texture[4][52] = 1;	green_platform_transparency_texture[4][53] = 1;	green_platform_transparency_texture[4][54] = 1;	green_platform_transparency_texture[4][55] = 1;	green_platform_transparency_texture[4][56] = 1;	green_platform_transparency_texture[4][57] = 1;	green_platform_transparency_texture[4][58] = 1;	green_platform_transparency_texture[4][59] = 1;	green_platform_transparency_texture[4][60] = 1;	green_platform_transparency_texture[4][61] = 1;	green_platform_transparency_texture[4][62] = 1;	green_platform_transparency_texture[4][63] = 1;	green_platform_transparency_texture[4][64] = 1;	green_platform_transparency_texture[4][65] = 1;	green_platform_transparency_texture[4][66] = 1;	green_platform_transparency_texture[4][67] = 1;	green_platform_transparency_texture[4][68] = 1;	green_platform_transparency_texture[4][69] = 1;	green_platform_transparency_texture[4][70] = 1;	green_platform_transparency_texture[4][71] = 1;	green_platform_transparency_texture[4][72] = 1;	green_platform_transparency_texture[4][73] = 1;	green_platform_transparency_texture[4][74] = 1;	green_platform_transparency_texture[4][75] = 1;	green_platform_transparency_texture[4][76] = 1;	green_platform_transparency_texture[4][77] = 1;	green_platform_transparency_texture[4][78] = 1;	green_platform_transparency_texture[4][79] = 1;	green_platform_transparency_texture[4][80] = 1;	green_platform_transparency_texture[4][81] = 1;	green_platform_transparency_texture[4][82] = 1;	green_platform_transparency_texture[4][83] = 1;	green_platform_transparency_texture[4][84] = 1;	green_platform_transparency_texture[4][85] = 1;	green_platform_transparency_texture[4][86] = 1;	green_platform_transparency_texture[4][87] = 1;	green_platform_transparency_texture[4][88] = 1;	green_platform_transparency_texture[4][89] = 1;	green_platform_transparency_texture[4][90] = 1;	green_platform_transparency_texture[4][91] = 1;	green_platform_transparency_texture[4][92] = 1;	green_platform_transparency_texture[4][93] = 1;	green_platform_transparency_texture[4][94] = 1;	green_platform_transparency_texture[4][95] = 1;	green_platform_transparency_texture[4][96] = 1;	green_platform_transparency_texture[4][97] = 1;	green_platform_transparency_texture[4][98] = 1;	green_platform_transparency_texture[4][99] = 1;	green_platform_transparency_texture[5][0] = 1;	green_platform_transparency_texture[5][1] = 1;	green_platform_transparency_texture[5][2] = 1;	green_platform_transparency_texture[5][3] = 1;	green_platform_transparency_texture[5][4] = 1;	green_platform_transparency_texture[5][5] = 1;	green_platform_transparency_texture[5][6] = 1;	green_platform_transparency_texture[5][7] = 1;	green_platform_transparency_texture[5][8] = 1;	green_platform_transparency_texture[5][9] = 1;	green_platform_transparency_texture[5][10] = 0;	green_platform_transparency_texture[5][11] = 0;	green_platform_transparency_texture[5][12] = 0;	green_platform_transparency_texture[5][13] = 0;	green_platform_transparency_texture[5][14] = 0;	green_platform_transparency_texture[5][15] = 0;	green_platform_transparency_texture[5][16] = 0;	green_platform_transparency_texture[5][17] = 0;	green_platform_transparency_texture[5][18] = 0;	green_platform_transparency_texture[5][19] = 0;	green_platform_transparency_texture[5][20] = 0;	green_platform_transparency_texture[5][21] = 0;	green_platform_transparency_texture[5][22] = 0;	green_platform_transparency_texture[5][23] = 0;	green_platform_transparency_texture[5][24] = 0;	green_platform_transparency_texture[5][25] = 0;	green_platform_transparency_texture[5][26] = 0;	green_platform_transparency_texture[5][27] = 0;	green_platform_transparency_texture[5][28] = 0;	green_platform_transparency_texture[5][29] = 0;	green_platform_transparency_texture[5][30] = 0;	green_platform_transparency_texture[5][31] = 0;	green_platform_transparency_texture[5][32] = 0;	green_platform_transparency_texture[5][33] = 0;	green_platform_transparency_texture[5][34] = 0;	green_platform_transparency_texture[5][35] = 0;	green_platform_transparency_texture[5][36] = 0;	green_platform_transparency_texture[5][37] = 0;	green_platform_transparency_texture[5][38] = 0;	green_platform_transparency_texture[5][39] = 0;	green_platform_transparency_texture[5][40] = 0;	green_platform_transparency_texture[5][41] = 0;	green_platform_transparency_texture[5][42] = 0;	green_platform_transparency_texture[5][43] = 0;	green_platform_transparency_texture[5][44] = 0;	green_platform_transparency_texture[5][45] = 0;	green_platform_transparency_texture[5][46] = 0;	green_platform_transparency_texture[5][47] = 0;	green_platform_transparency_texture[5][48] = 0;	green_platform_transparency_texture[5][49] = 0;	green_platform_transparency_texture[5][50] = 0;	green_platform_transparency_texture[5][51] = 0;	green_platform_transparency_texture[5][52] = 0;	green_platform_transparency_texture[5][53] = 0;	green_platform_transparency_texture[5][54] = 0;	green_platform_transparency_texture[5][55] = 0;	green_platform_transparency_texture[5][56] = 0;	green_platform_transparency_texture[5][57] = 0;	green_platform_transparency_texture[5][58] = 0;	green_platform_transparency_texture[5][59] = 0;	green_platform_transparency_texture[5][60] = 0;	green_platform_transparency_texture[5][61] = 0;	green_platform_transparency_texture[5][62] = 0;	green_platform_transparency_texture[5][63] = 0;	green_platform_transparency_texture[5][64] = 0;	green_platform_transparency_texture[5][65] = 0;	green_platform_transparency_texture[5][66] = 0;	green_platform_transparency_texture[5][67] = 0;	green_platform_transparency_texture[5][68] = 0;	green_platform_transparency_texture[5][69] = 0;	green_platform_transparency_texture[5][70] = 0;	green_platform_transparency_texture[5][71] = 0;	green_platform_transparency_texture[5][72] = 0;	green_platform_transparency_texture[5][73] = 0;	green_platform_transparency_texture[5][74] = 0;	green_platform_transparency_texture[5][75] = 0;	green_platform_transparency_texture[5][76] = 0;	green_platform_transparency_texture[5][77] = 0;	green_platform_transparency_texture[5][78] = 0;	green_platform_transparency_texture[5][79] = 0;	green_platform_transparency_texture[5][80] = 0;	green_platform_transparency_texture[5][81] = 0;	green_platform_transparency_texture[5][82] = 0;	green_platform_transparency_texture[5][83] = 0;	green_platform_transparency_texture[5][84] = 0;	green_platform_transparency_texture[5][85] = 0;	green_platform_transparency_texture[5][86] = 0;	green_platform_transparency_texture[5][87] = 0;	green_platform_transparency_texture[5][88] = 0;	green_platform_transparency_texture[5][89] = 0;	green_platform_transparency_texture[5][90] = 1;	green_platform_transparency_texture[5][91] = 1;	green_platform_transparency_texture[5][92] = 1;	green_platform_transparency_texture[5][93] = 1;	green_platform_transparency_texture[5][94] = 1;	green_platform_transparency_texture[5][95] = 1;	green_platform_transparency_texture[5][96] = 1;	green_platform_transparency_texture[5][97] = 1;	green_platform_transparency_texture[5][98] = 1;	green_platform_transparency_texture[5][99] = 1;	green_platform_transparency_texture[6][0] = 1;	green_platform_transparency_texture[6][1] = 1;	green_platform_transparency_texture[6][2] = 1;	green_platform_transparency_texture[6][3] = 1;	green_platform_transparency_texture[6][4] = 1;	green_platform_transparency_texture[6][5] = 1;	green_platform_transparency_texture[6][6] = 1;	green_platform_transparency_texture[6][7] = 1;	green_platform_transparency_texture[6][8] = 1;	green_platform_transparency_texture[6][9] = 1;	green_platform_transparency_texture[6][10] = 0;	green_platform_transparency_texture[6][11] = 0;	green_platform_transparency_texture[6][12] = 0;	green_platform_transparency_texture[6][13] = 0;	green_platform_transparency_texture[6][14] = 0;	green_platform_transparency_texture[6][15] = 0;	green_platform_transparency_texture[6][16] = 0;	green_platform_transparency_texture[6][17] = 0;	green_platform_transparency_texture[6][18] = 0;	green_platform_transparency_texture[6][19] = 0;	green_platform_transparency_texture[6][20] = 0;	green_platform_transparency_texture[6][21] = 0;	green_platform_transparency_texture[6][22] = 0;	green_platform_transparency_texture[6][23] = 0;	green_platform_transparency_texture[6][24] = 0;	green_platform_transparency_texture[6][25] = 0;	green_platform_transparency_texture[6][26] = 0;	green_platform_transparency_texture[6][27] = 0;	green_platform_transparency_texture[6][28] = 0;	green_platform_transparency_texture[6][29] = 0;	green_platform_transparency_texture[6][30] = 0;	green_platform_transparency_texture[6][31] = 0;	green_platform_transparency_texture[6][32] = 0;	green_platform_transparency_texture[6][33] = 0;	green_platform_transparency_texture[6][34] = 0;	green_platform_transparency_texture[6][35] = 0;	green_platform_transparency_texture[6][36] = 0;	green_platform_transparency_texture[6][37] = 0;	green_platform_transparency_texture[6][38] = 0;	green_platform_transparency_texture[6][39] = 0;	green_platform_transparency_texture[6][40] = 0;	green_platform_transparency_texture[6][41] = 0;	green_platform_transparency_texture[6][42] = 0;	green_platform_transparency_texture[6][43] = 0;	green_platform_transparency_texture[6][44] = 0;	green_platform_transparency_texture[6][45] = 0;	green_platform_transparency_texture[6][46] = 0;	green_platform_transparency_texture[6][47] = 0;	green_platform_transparency_texture[6][48] = 0;	green_platform_transparency_texture[6][49] = 0;	green_platform_transparency_texture[6][50] = 0;	green_platform_transparency_texture[6][51] = 0;	green_platform_transparency_texture[6][52] = 0;	green_platform_transparency_texture[6][53] = 0;	green_platform_transparency_texture[6][54] = 0;	green_platform_transparency_texture[6][55] = 0;	green_platform_transparency_texture[6][56] = 0;	green_platform_transparency_texture[6][57] = 0;	green_platform_transparency_texture[6][58] = 0;	green_platform_transparency_texture[6][59] = 0;	green_platform_transparency_texture[6][60] = 0;	green_platform_transparency_texture[6][61] = 0;	green_platform_transparency_texture[6][62] = 0;	green_platform_transparency_texture[6][63] = 0;	green_platform_transparency_texture[6][64] = 0;	green_platform_transparency_texture[6][65] = 0;	green_platform_transparency_texture[6][66] = 0;	green_platform_transparency_texture[6][67] = 0;	green_platform_transparency_texture[6][68] = 0;	green_platform_transparency_texture[6][69] = 0;	green_platform_transparency_texture[6][70] = 0;	green_platform_transparency_texture[6][71] = 0;	green_platform_transparency_texture[6][72] = 0;	green_platform_transparency_texture[6][73] = 0;	green_platform_transparency_texture[6][74] = 0;	green_platform_transparency_texture[6][75] = 0;	green_platform_transparency_texture[6][76] = 0;	green_platform_transparency_texture[6][77] = 0;	green_platform_transparency_texture[6][78] = 0;	green_platform_transparency_texture[6][79] = 0;	green_platform_transparency_texture[6][80] = 0;	green_platform_transparency_texture[6][81] = 0;	green_platform_transparency_texture[6][82] = 0;	green_platform_transparency_texture[6][83] = 0;	green_platform_transparency_texture[6][84] = 0;	green_platform_transparency_texture[6][85] = 0;	green_platform_transparency_texture[6][86] = 0;	green_platform_transparency_texture[6][87] = 0;	green_platform_transparency_texture[6][88] = 0;	green_platform_transparency_texture[6][89] = 0;	green_platform_transparency_texture[6][90] = 1;	green_platform_transparency_texture[6][91] = 1;	green_platform_transparency_texture[6][92] = 1;	green_platform_transparency_texture[6][93] = 1;	green_platform_transparency_texture[6][94] = 1;	green_platform_transparency_texture[6][95] = 1;	green_platform_transparency_texture[6][96] = 1;	green_platform_transparency_texture[6][97] = 1;	green_platform_transparency_texture[6][98] = 1;	green_platform_transparency_texture[6][99] = 1;	green_platform_transparency_texture[7][0] = 1;	green_platform_transparency_texture[7][1] = 1;	green_platform_transparency_texture[7][2] = 1;	green_platform_transparency_texture[7][3] = 1;	green_platform_transparency_texture[7][4] = 1;	green_platform_transparency_texture[7][5] = 1;	green_platform_transparency_texture[7][6] = 1;	green_platform_transparency_texture[7][7] = 1;	green_platform_transparency_texture[7][8] = 1;	green_platform_transparency_texture[7][9] = 1;	green_platform_transparency_texture[7][10] = 0;	green_platform_transparency_texture[7][11] = 0;	green_platform_transparency_texture[7][12] = 0;	green_platform_transparency_texture[7][13] = 0;	green_platform_transparency_texture[7][14] = 0;	green_platform_transparency_texture[7][15] = 0;	green_platform_transparency_texture[7][16] = 0;	green_platform_transparency_texture[7][17] = 0;	green_platform_transparency_texture[7][18] = 0;	green_platform_transparency_texture[7][19] = 0;	green_platform_transparency_texture[7][20] = 0;	green_platform_transparency_texture[7][21] = 0;	green_platform_transparency_texture[7][22] = 0;	green_platform_transparency_texture[7][23] = 0;	green_platform_transparency_texture[7][24] = 0;	green_platform_transparency_texture[7][25] = 0;	green_platform_transparency_texture[7][26] = 0;	green_platform_transparency_texture[7][27] = 0;	green_platform_transparency_texture[7][28] = 0;	green_platform_transparency_texture[7][29] = 0;	green_platform_transparency_texture[7][30] = 0;	green_platform_transparency_texture[7][31] = 0;	green_platform_transparency_texture[7][32] = 0;	green_platform_transparency_texture[7][33] = 0;	green_platform_transparency_texture[7][34] = 0;	green_platform_transparency_texture[7][35] = 0;	green_platform_transparency_texture[7][36] = 0;	green_platform_transparency_texture[7][37] = 0;	green_platform_transparency_texture[7][38] = 0;	green_platform_transparency_texture[7][39] = 0;	green_platform_transparency_texture[7][40] = 0;	green_platform_transparency_texture[7][41] = 0;	green_platform_transparency_texture[7][42] = 0;	green_platform_transparency_texture[7][43] = 0;	green_platform_transparency_texture[7][44] = 0;	green_platform_transparency_texture[7][45] = 0;	green_platform_transparency_texture[7][46] = 0;	green_platform_transparency_texture[7][47] = 0;	green_platform_transparency_texture[7][48] = 0;	green_platform_transparency_texture[7][49] = 0;	green_platform_transparency_texture[7][50] = 0;	green_platform_transparency_texture[7][51] = 0;	green_platform_transparency_texture[7][52] = 0;	green_platform_transparency_texture[7][53] = 0;	green_platform_transparency_texture[7][54] = 0;	green_platform_transparency_texture[7][55] = 0;	green_platform_transparency_texture[7][56] = 0;	green_platform_transparency_texture[7][57] = 0;	green_platform_transparency_texture[7][58] = 0;	green_platform_transparency_texture[7][59] = 0;	green_platform_transparency_texture[7][60] = 0;	green_platform_transparency_texture[7][61] = 0;	green_platform_transparency_texture[7][62] = 0;	green_platform_transparency_texture[7][63] = 0;	green_platform_transparency_texture[7][64] = 0;	green_platform_transparency_texture[7][65] = 0;	green_platform_transparency_texture[7][66] = 0;	green_platform_transparency_texture[7][67] = 0;	green_platform_transparency_texture[7][68] = 0;	green_platform_transparency_texture[7][69] = 0;	green_platform_transparency_texture[7][70] = 0;	green_platform_transparency_texture[7][71] = 0;	green_platform_transparency_texture[7][72] = 0;	green_platform_transparency_texture[7][73] = 0;	green_platform_transparency_texture[7][74] = 0;	green_platform_transparency_texture[7][75] = 0;	green_platform_transparency_texture[7][76] = 0;	green_platform_transparency_texture[7][77] = 0;	green_platform_transparency_texture[7][78] = 0;	green_platform_transparency_texture[7][79] = 0;	green_platform_transparency_texture[7][80] = 0;	green_platform_transparency_texture[7][81] = 0;	green_platform_transparency_texture[7][82] = 0;	green_platform_transparency_texture[7][83] = 0;	green_platform_transparency_texture[7][84] = 0;	green_platform_transparency_texture[7][85] = 0;	green_platform_transparency_texture[7][86] = 0;	green_platform_transparency_texture[7][87] = 0;	green_platform_transparency_texture[7][88] = 0;	green_platform_transparency_texture[7][89] = 0;	green_platform_transparency_texture[7][90] = 1;	green_platform_transparency_texture[7][91] = 1;	green_platform_transparency_texture[7][92] = 1;	green_platform_transparency_texture[7][93] = 1;	green_platform_transparency_texture[7][94] = 1;	green_platform_transparency_texture[7][95] = 1;	green_platform_transparency_texture[7][96] = 1;	green_platform_transparency_texture[7][97] = 1;	green_platform_transparency_texture[7][98] = 1;	green_platform_transparency_texture[7][99] = 1;	green_platform_transparency_texture[8][0] = 1;	green_platform_transparency_texture[8][1] = 1;	green_platform_transparency_texture[8][2] = 1;	green_platform_transparency_texture[8][3] = 1;	green_platform_transparency_texture[8][4] = 1;	green_platform_transparency_texture[8][5] = 1;	green_platform_transparency_texture[8][6] = 1;	green_platform_transparency_texture[8][7] = 1;	green_platform_transparency_texture[8][8] = 1;	green_platform_transparency_texture[8][9] = 1;	green_platform_transparency_texture[8][10] = 0;	green_platform_transparency_texture[8][11] = 0;	green_platform_transparency_texture[8][12] = 0;	green_platform_transparency_texture[8][13] = 0;	green_platform_transparency_texture[8][14] = 0;	green_platform_transparency_texture[8][15] = 0;	green_platform_transparency_texture[8][16] = 0;	green_platform_transparency_texture[8][17] = 0;	green_platform_transparency_texture[8][18] = 0;	green_platform_transparency_texture[8][19] = 0;	green_platform_transparency_texture[8][20] = 0;	green_platform_transparency_texture[8][21] = 0;	green_platform_transparency_texture[8][22] = 0;	green_platform_transparency_texture[8][23] = 0;	green_platform_transparency_texture[8][24] = 0;	green_platform_transparency_texture[8][25] = 0;	green_platform_transparency_texture[8][26] = 0;	green_platform_transparency_texture[8][27] = 0;	green_platform_transparency_texture[8][28] = 0;	green_platform_transparency_texture[8][29] = 0;	green_platform_transparency_texture[8][30] = 0;	green_platform_transparency_texture[8][31] = 0;	green_platform_transparency_texture[8][32] = 0;	green_platform_transparency_texture[8][33] = 0;	green_platform_transparency_texture[8][34] = 0;	green_platform_transparency_texture[8][35] = 0;	green_platform_transparency_texture[8][36] = 0;	green_platform_transparency_texture[8][37] = 0;	green_platform_transparency_texture[8][38] = 0;	green_platform_transparency_texture[8][39] = 0;	green_platform_transparency_texture[8][40] = 0;	green_platform_transparency_texture[8][41] = 0;	green_platform_transparency_texture[8][42] = 0;	green_platform_transparency_texture[8][43] = 0;	green_platform_transparency_texture[8][44] = 0;	green_platform_transparency_texture[8][45] = 0;	green_platform_transparency_texture[8][46] = 0;	green_platform_transparency_texture[8][47] = 0;	green_platform_transparency_texture[8][48] = 0;	green_platform_transparency_texture[8][49] = 0;	green_platform_transparency_texture[8][50] = 0;	green_platform_transparency_texture[8][51] = 0;	green_platform_transparency_texture[8][52] = 0;	green_platform_transparency_texture[8][53] = 0;	green_platform_transparency_texture[8][54] = 0;	green_platform_transparency_texture[8][55] = 0;	green_platform_transparency_texture[8][56] = 0;	green_platform_transparency_texture[8][57] = 0;	green_platform_transparency_texture[8][58] = 0;	green_platform_transparency_texture[8][59] = 0;	green_platform_transparency_texture[8][60] = 0;	green_platform_transparency_texture[8][61] = 0;	green_platform_transparency_texture[8][62] = 0;	green_platform_transparency_texture[8][63] = 0;	green_platform_transparency_texture[8][64] = 0;	green_platform_transparency_texture[8][65] = 0;	green_platform_transparency_texture[8][66] = 0;	green_platform_transparency_texture[8][67] = 0;	green_platform_transparency_texture[8][68] = 0;	green_platform_transparency_texture[8][69] = 0;	green_platform_transparency_texture[8][70] = 0;	green_platform_transparency_texture[8][71] = 0;	green_platform_transparency_texture[8][72] = 0;	green_platform_transparency_texture[8][73] = 0;	green_platform_transparency_texture[8][74] = 0;	green_platform_transparency_texture[8][75] = 0;	green_platform_transparency_texture[8][76] = 0;	green_platform_transparency_texture[8][77] = 0;	green_platform_transparency_texture[8][78] = 0;	green_platform_transparency_texture[8][79] = 0;	green_platform_transparency_texture[8][80] = 0;	green_platform_transparency_texture[8][81] = 0;	green_platform_transparency_texture[8][82] = 0;	green_platform_transparency_texture[8][83] = 0;	green_platform_transparency_texture[8][84] = 0;	green_platform_transparency_texture[8][85] = 0;	green_platform_transparency_texture[8][86] = 0;	green_platform_transparency_texture[8][87] = 0;	green_platform_transparency_texture[8][88] = 0;	green_platform_transparency_texture[8][89] = 0;	green_platform_transparency_texture[8][90] = 1;	green_platform_transparency_texture[8][91] = 1;	green_platform_transparency_texture[8][92] = 1;	green_platform_transparency_texture[8][93] = 1;	green_platform_transparency_texture[8][94] = 1;	green_platform_transparency_texture[8][95] = 1;	green_platform_transparency_texture[8][96] = 1;	green_platform_transparency_texture[8][97] = 1;	green_platform_transparency_texture[8][98] = 1;	green_platform_transparency_texture[8][99] = 1;	green_platform_transparency_texture[9][0] = 1;	green_platform_transparency_texture[9][1] = 1;	green_platform_transparency_texture[9][2] = 1;	green_platform_transparency_texture[9][3] = 1;	green_platform_transparency_texture[9][4] = 1;	green_platform_transparency_texture[9][5] = 1;	green_platform_transparency_texture[9][6] = 1;	green_platform_transparency_texture[9][7] = 1;	green_platform_transparency_texture[9][8] = 1;	green_platform_transparency_texture[9][9] = 1;	green_platform_transparency_texture[9][10] = 0;	green_platform_transparency_texture[9][11] = 0;	green_platform_transparency_texture[9][12] = 0;	green_platform_transparency_texture[9][13] = 0;	green_platform_transparency_texture[9][14] = 0;	green_platform_transparency_texture[9][15] = 0;	green_platform_transparency_texture[9][16] = 0;	green_platform_transparency_texture[9][17] = 0;	green_platform_transparency_texture[9][18] = 0;	green_platform_transparency_texture[9][19] = 0;	green_platform_transparency_texture[9][20] = 0;	green_platform_transparency_texture[9][21] = 0;	green_platform_transparency_texture[9][22] = 0;	green_platform_transparency_texture[9][23] = 0;	green_platform_transparency_texture[9][24] = 0;	green_platform_transparency_texture[9][25] = 0;	green_platform_transparency_texture[9][26] = 0;	green_platform_transparency_texture[9][27] = 0;	green_platform_transparency_texture[9][28] = 0;	green_platform_transparency_texture[9][29] = 0;	green_platform_transparency_texture[9][30] = 0;	green_platform_transparency_texture[9][31] = 0;	green_platform_transparency_texture[9][32] = 0;	green_platform_transparency_texture[9][33] = 0;	green_platform_transparency_texture[9][34] = 0;	green_platform_transparency_texture[9][35] = 0;	green_platform_transparency_texture[9][36] = 0;	green_platform_transparency_texture[9][37] = 0;	green_platform_transparency_texture[9][38] = 0;	green_platform_transparency_texture[9][39] = 0;	green_platform_transparency_texture[9][40] = 0;	green_platform_transparency_texture[9][41] = 0;	green_platform_transparency_texture[9][42] = 0;	green_platform_transparency_texture[9][43] = 0;	green_platform_transparency_texture[9][44] = 0;	green_platform_transparency_texture[9][45] = 0;	green_platform_transparency_texture[9][46] = 0;	green_platform_transparency_texture[9][47] = 0;	green_platform_transparency_texture[9][48] = 0;	green_platform_transparency_texture[9][49] = 0;	green_platform_transparency_texture[9][50] = 0;	green_platform_transparency_texture[9][51] = 0;	green_platform_transparency_texture[9][52] = 0;	green_platform_transparency_texture[9][53] = 0;	green_platform_transparency_texture[9][54] = 0;	green_platform_transparency_texture[9][55] = 0;	green_platform_transparency_texture[9][56] = 0;	green_platform_transparency_texture[9][57] = 0;	green_platform_transparency_texture[9][58] = 0;	green_platform_transparency_texture[9][59] = 0;	green_platform_transparency_texture[9][60] = 0;	green_platform_transparency_texture[9][61] = 0;	green_platform_transparency_texture[9][62] = 0;	green_platform_transparency_texture[9][63] = 0;	green_platform_transparency_texture[9][64] = 0;	green_platform_transparency_texture[9][65] = 0;	green_platform_transparency_texture[9][66] = 0;	green_platform_transparency_texture[9][67] = 0;	green_platform_transparency_texture[9][68] = 0;	green_platform_transparency_texture[9][69] = 0;	green_platform_transparency_texture[9][70] = 0;	green_platform_transparency_texture[9][71] = 0;	green_platform_transparency_texture[9][72] = 0;	green_platform_transparency_texture[9][73] = 0;	green_platform_transparency_texture[9][74] = 0;	green_platform_transparency_texture[9][75] = 0;	green_platform_transparency_texture[9][76] = 0;	green_platform_transparency_texture[9][77] = 0;	green_platform_transparency_texture[9][78] = 0;	green_platform_transparency_texture[9][79] = 0;	green_platform_transparency_texture[9][80] = 0;	green_platform_transparency_texture[9][81] = 0;	green_platform_transparency_texture[9][82] = 0;	green_platform_transparency_texture[9][83] = 0;	green_platform_transparency_texture[9][84] = 0;	green_platform_transparency_texture[9][85] = 0;	green_platform_transparency_texture[9][86] = 0;	green_platform_transparency_texture[9][87] = 0;	green_platform_transparency_texture[9][88] = 0;	green_platform_transparency_texture[9][89] = 0;	green_platform_transparency_texture[9][90] = 1;	green_platform_transparency_texture[9][91] = 1;	green_platform_transparency_texture[9][92] = 1;	green_platform_transparency_texture[9][93] = 1;	green_platform_transparency_texture[9][94] = 1;	green_platform_transparency_texture[9][95] = 1;	green_platform_transparency_texture[9][96] = 1;	green_platform_transparency_texture[9][97] = 1;	green_platform_transparency_texture[9][98] = 1;	green_platform_transparency_texture[9][99] = 1;	green_platform_transparency_texture[10][0] = 1;	green_platform_transparency_texture[10][1] = 1;	green_platform_transparency_texture[10][2] = 1;	green_platform_transparency_texture[10][3] = 1;	green_platform_transparency_texture[10][4] = 1;	green_platform_transparency_texture[10][5] = 0;	green_platform_transparency_texture[10][6] = 0;	green_platform_transparency_texture[10][7] = 0;	green_platform_transparency_texture[10][8] = 0;	green_platform_transparency_texture[10][9] = 0;	green_platform_transparency_texture[10][10] = 0;	green_platform_transparency_texture[10][11] = 0;	green_platform_transparency_texture[10][12] = 0;	green_platform_transparency_texture[10][13] = 0;	green_platform_transparency_texture[10][14] = 0;	green_platform_transparency_texture[10][15] = 0;	green_platform_transparency_texture[10][16] = 0;	green_platform_transparency_texture[10][17] = 0;	green_platform_transparency_texture[10][18] = 0;	green_platform_transparency_texture[10][19] = 0;	green_platform_transparency_texture[10][20] = 0;	green_platform_transparency_texture[10][21] = 0;	green_platform_transparency_texture[10][22] = 0;	green_platform_transparency_texture[10][23] = 0;	green_platform_transparency_texture[10][24] = 0;	green_platform_transparency_texture[10][25] = 0;	green_platform_transparency_texture[10][26] = 0;	green_platform_transparency_texture[10][27] = 0;	green_platform_transparency_texture[10][28] = 0;	green_platform_transparency_texture[10][29] = 0;	green_platform_transparency_texture[10][30] = 0;	green_platform_transparency_texture[10][31] = 0;	green_platform_transparency_texture[10][32] = 0;	green_platform_transparency_texture[10][33] = 0;	green_platform_transparency_texture[10][34] = 0;	green_platform_transparency_texture[10][35] = 0;	green_platform_transparency_texture[10][36] = 0;	green_platform_transparency_texture[10][37] = 0;	green_platform_transparency_texture[10][38] = 0;	green_platform_transparency_texture[10][39] = 0;	green_platform_transparency_texture[10][40] = 0;	green_platform_transparency_texture[10][41] = 0;	green_platform_transparency_texture[10][42] = 0;	green_platform_transparency_texture[10][43] = 0;	green_platform_transparency_texture[10][44] = 0;	green_platform_transparency_texture[10][45] = 0;	green_platform_transparency_texture[10][46] = 0;	green_platform_transparency_texture[10][47] = 0;	green_platform_transparency_texture[10][48] = 0;	green_platform_transparency_texture[10][49] = 0;	green_platform_transparency_texture[10][50] = 0;	green_platform_transparency_texture[10][51] = 0;	green_platform_transparency_texture[10][52] = 0;	green_platform_transparency_texture[10][53] = 0;	green_platform_transparency_texture[10][54] = 0;	green_platform_transparency_texture[10][55] = 0;	green_platform_transparency_texture[10][56] = 0;	green_platform_transparency_texture[10][57] = 0;	green_platform_transparency_texture[10][58] = 0;	green_platform_transparency_texture[10][59] = 0;	green_platform_transparency_texture[10][60] = 0;	green_platform_transparency_texture[10][61] = 0;	green_platform_transparency_texture[10][62] = 0;	green_platform_transparency_texture[10][63] = 0;	green_platform_transparency_texture[10][64] = 0;	green_platform_transparency_texture[10][65] = 0;	green_platform_transparency_texture[10][66] = 0;	green_platform_transparency_texture[10][67] = 0;	green_platform_transparency_texture[10][68] = 0;	green_platform_transparency_texture[10][69] = 0;	green_platform_transparency_texture[10][70] = 0;	green_platform_transparency_texture[10][71] = 0;	green_platform_transparency_texture[10][72] = 0;	green_platform_transparency_texture[10][73] = 0;	green_platform_transparency_texture[10][74] = 0;	green_platform_transparency_texture[10][75] = 0;	green_platform_transparency_texture[10][76] = 0;	green_platform_transparency_texture[10][77] = 0;	green_platform_transparency_texture[10][78] = 0;	green_platform_transparency_texture[10][79] = 0;	green_platform_transparency_texture[10][80] = 0;	green_platform_transparency_texture[10][81] = 0;	green_platform_transparency_texture[10][82] = 0;	green_platform_transparency_texture[10][83] = 0;	green_platform_transparency_texture[10][84] = 0;	green_platform_transparency_texture[10][85] = 0;	green_platform_transparency_texture[10][86] = 0;	green_platform_transparency_texture[10][87] = 0;	green_platform_transparency_texture[10][88] = 0;	green_platform_transparency_texture[10][89] = 0;	green_platform_transparency_texture[10][90] = 0;	green_platform_transparency_texture[10][91] = 0;	green_platform_transparency_texture[10][92] = 0;	green_platform_transparency_texture[10][93] = 0;	green_platform_transparency_texture[10][94] = 0;	green_platform_transparency_texture[10][95] = 1;	green_platform_transparency_texture[10][96] = 1;	green_platform_transparency_texture[10][97] = 1;	green_platform_transparency_texture[10][98] = 1;	green_platform_transparency_texture[10][99] = 1;	green_platform_transparency_texture[11][0] = 1;	green_platform_transparency_texture[11][1] = 1;	green_platform_transparency_texture[11][2] = 1;	green_platform_transparency_texture[11][3] = 1;	green_platform_transparency_texture[11][4] = 1;	green_platform_transparency_texture[11][5] = 0;	green_platform_transparency_texture[11][6] = 0;	green_platform_transparency_texture[11][7] = 0;	green_platform_transparency_texture[11][8] = 0;	green_platform_transparency_texture[11][9] = 0;	green_platform_transparency_texture[11][10] = 0;	green_platform_transparency_texture[11][11] = 0;	green_platform_transparency_texture[11][12] = 0;	green_platform_transparency_texture[11][13] = 0;	green_platform_transparency_texture[11][14] = 0;	green_platform_transparency_texture[11][15] = 0;	green_platform_transparency_texture[11][16] = 0;	green_platform_transparency_texture[11][17] = 0;	green_platform_transparency_texture[11][18] = 0;	green_platform_transparency_texture[11][19] = 0;	green_platform_transparency_texture[11][20] = 0;	green_platform_transparency_texture[11][21] = 0;	green_platform_transparency_texture[11][22] = 0;	green_platform_transparency_texture[11][23] = 0;	green_platform_transparency_texture[11][24] = 0;	green_platform_transparency_texture[11][25] = 0;	green_platform_transparency_texture[11][26] = 0;	green_platform_transparency_texture[11][27] = 0;	green_platform_transparency_texture[11][28] = 0;	green_platform_transparency_texture[11][29] = 0;	green_platform_transparency_texture[11][30] = 0;	green_platform_transparency_texture[11][31] = 0;	green_platform_transparency_texture[11][32] = 0;	green_platform_transparency_texture[11][33] = 0;	green_platform_transparency_texture[11][34] = 0;	green_platform_transparency_texture[11][35] = 0;	green_platform_transparency_texture[11][36] = 0;	green_platform_transparency_texture[11][37] = 0;	green_platform_transparency_texture[11][38] = 0;	green_platform_transparency_texture[11][39] = 0;	green_platform_transparency_texture[11][40] = 0;	green_platform_transparency_texture[11][41] = 0;	green_platform_transparency_texture[11][42] = 0;	green_platform_transparency_texture[11][43] = 0;	green_platform_transparency_texture[11][44] = 0;	green_platform_transparency_texture[11][45] = 0;	green_platform_transparency_texture[11][46] = 0;	green_platform_transparency_texture[11][47] = 0;	green_platform_transparency_texture[11][48] = 0;	green_platform_transparency_texture[11][49] = 0;	green_platform_transparency_texture[11][50] = 0;	green_platform_transparency_texture[11][51] = 0;	green_platform_transparency_texture[11][52] = 0;	green_platform_transparency_texture[11][53] = 0;	green_platform_transparency_texture[11][54] = 0;	green_platform_transparency_texture[11][55] = 0;	green_platform_transparency_texture[11][56] = 0;	green_platform_transparency_texture[11][57] = 0;	green_platform_transparency_texture[11][58] = 0;	green_platform_transparency_texture[11][59] = 0;	green_platform_transparency_texture[11][60] = 0;	green_platform_transparency_texture[11][61] = 0;	green_platform_transparency_texture[11][62] = 0;	green_platform_transparency_texture[11][63] = 0;	green_platform_transparency_texture[11][64] = 0;	green_platform_transparency_texture[11][65] = 0;	green_platform_transparency_texture[11][66] = 0;	green_platform_transparency_texture[11][67] = 0;	green_platform_transparency_texture[11][68] = 0;	green_platform_transparency_texture[11][69] = 0;	green_platform_transparency_texture[11][70] = 0;	green_platform_transparency_texture[11][71] = 0;	green_platform_transparency_texture[11][72] = 0;	green_platform_transparency_texture[11][73] = 0;	green_platform_transparency_texture[11][74] = 0;	green_platform_transparency_texture[11][75] = 0;	green_platform_transparency_texture[11][76] = 0;	green_platform_transparency_texture[11][77] = 0;	green_platform_transparency_texture[11][78] = 0;	green_platform_transparency_texture[11][79] = 0;	green_platform_transparency_texture[11][80] = 0;	green_platform_transparency_texture[11][81] = 0;	green_platform_transparency_texture[11][82] = 0;	green_platform_transparency_texture[11][83] = 0;	green_platform_transparency_texture[11][84] = 0;	green_platform_transparency_texture[11][85] = 0;	green_platform_transparency_texture[11][86] = 0;	green_platform_transparency_texture[11][87] = 0;	green_platform_transparency_texture[11][88] = 0;	green_platform_transparency_texture[11][89] = 0;	green_platform_transparency_texture[11][90] = 0;	green_platform_transparency_texture[11][91] = 0;	green_platform_transparency_texture[11][92] = 0;	green_platform_transparency_texture[11][93] = 0;	green_platform_transparency_texture[11][94] = 0;	green_platform_transparency_texture[11][95] = 1;	green_platform_transparency_texture[11][96] = 1;	green_platform_transparency_texture[11][97] = 1;	green_platform_transparency_texture[11][98] = 1;	green_platform_transparency_texture[11][99] = 1;	green_platform_transparency_texture[12][0] = 1;	green_platform_transparency_texture[12][1] = 1;	green_platform_transparency_texture[12][2] = 1;	green_platform_transparency_texture[12][3] = 1;	green_platform_transparency_texture[12][4] = 1;	green_platform_transparency_texture[12][5] = 0;	green_platform_transparency_texture[12][6] = 0;	green_platform_transparency_texture[12][7] = 0;	green_platform_transparency_texture[12][8] = 0;	green_platform_transparency_texture[12][9] = 0;	green_platform_transparency_texture[12][10] = 0;	green_platform_transparency_texture[12][11] = 0;	green_platform_transparency_texture[12][12] = 0;	green_platform_transparency_texture[12][13] = 0;	green_platform_transparency_texture[12][14] = 0;	green_platform_transparency_texture[12][15] = 0;	green_platform_transparency_texture[12][16] = 0;	green_platform_transparency_texture[12][17] = 0;	green_platform_transparency_texture[12][18] = 0;	green_platform_transparency_texture[12][19] = 0;	green_platform_transparency_texture[12][20] = 0;	green_platform_transparency_texture[12][21] = 0;	green_platform_transparency_texture[12][22] = 0;	green_platform_transparency_texture[12][23] = 0;	green_platform_transparency_texture[12][24] = 0;	green_platform_transparency_texture[12][25] = 0;	green_platform_transparency_texture[12][26] = 0;	green_platform_transparency_texture[12][27] = 0;	green_platform_transparency_texture[12][28] = 0;	green_platform_transparency_texture[12][29] = 0;	green_platform_transparency_texture[12][30] = 0;	green_platform_transparency_texture[12][31] = 0;	green_platform_transparency_texture[12][32] = 0;	green_platform_transparency_texture[12][33] = 0;	green_platform_transparency_texture[12][34] = 0;	green_platform_transparency_texture[12][35] = 0;	green_platform_transparency_texture[12][36] = 0;	green_platform_transparency_texture[12][37] = 0;	green_platform_transparency_texture[12][38] = 0;	green_platform_transparency_texture[12][39] = 0;	green_platform_transparency_texture[12][40] = 0;	green_platform_transparency_texture[12][41] = 0;	green_platform_transparency_texture[12][42] = 0;	green_platform_transparency_texture[12][43] = 0;	green_platform_transparency_texture[12][44] = 0;	green_platform_transparency_texture[12][45] = 0;	green_platform_transparency_texture[12][46] = 0;	green_platform_transparency_texture[12][47] = 0;	green_platform_transparency_texture[12][48] = 0;	green_platform_transparency_texture[12][49] = 0;	green_platform_transparency_texture[12][50] = 0;	green_platform_transparency_texture[12][51] = 0;	green_platform_transparency_texture[12][52] = 0;	green_platform_transparency_texture[12][53] = 0;	green_platform_transparency_texture[12][54] = 0;	green_platform_transparency_texture[12][55] = 0;	green_platform_transparency_texture[12][56] = 0;	green_platform_transparency_texture[12][57] = 0;	green_platform_transparency_texture[12][58] = 0;	green_platform_transparency_texture[12][59] = 0;	green_platform_transparency_texture[12][60] = 0;	green_platform_transparency_texture[12][61] = 0;	green_platform_transparency_texture[12][62] = 0;	green_platform_transparency_texture[12][63] = 0;	green_platform_transparency_texture[12][64] = 0;	green_platform_transparency_texture[12][65] = 0;	green_platform_transparency_texture[12][66] = 0;	green_platform_transparency_texture[12][67] = 0;	green_platform_transparency_texture[12][68] = 0;	green_platform_transparency_texture[12][69] = 0;	green_platform_transparency_texture[12][70] = 0;	green_platform_transparency_texture[12][71] = 0;	green_platform_transparency_texture[12][72] = 0;	green_platform_transparency_texture[12][73] = 0;	green_platform_transparency_texture[12][74] = 0;	green_platform_transparency_texture[12][75] = 0;	green_platform_transparency_texture[12][76] = 0;	green_platform_transparency_texture[12][77] = 0;	green_platform_transparency_texture[12][78] = 0;	green_platform_transparency_texture[12][79] = 0;	green_platform_transparency_texture[12][80] = 0;	green_platform_transparency_texture[12][81] = 0;	green_platform_transparency_texture[12][82] = 0;	green_platform_transparency_texture[12][83] = 0;	green_platform_transparency_texture[12][84] = 0;	green_platform_transparency_texture[12][85] = 0;	green_platform_transparency_texture[12][86] = 0;	green_platform_transparency_texture[12][87] = 0;	green_platform_transparency_texture[12][88] = 0;	green_platform_transparency_texture[12][89] = 0;	green_platform_transparency_texture[12][90] = 0;	green_platform_transparency_texture[12][91] = 0;	green_platform_transparency_texture[12][92] = 0;	green_platform_transparency_texture[12][93] = 0;	green_platform_transparency_texture[12][94] = 0;	green_platform_transparency_texture[12][95] = 1;	green_platform_transparency_texture[12][96] = 1;	green_platform_transparency_texture[12][97] = 1;	green_platform_transparency_texture[12][98] = 1;	green_platform_transparency_texture[12][99] = 1;	green_platform_transparency_texture[13][0] = 1;	green_platform_transparency_texture[13][1] = 1;	green_platform_transparency_texture[13][2] = 1;	green_platform_transparency_texture[13][3] = 1;	green_platform_transparency_texture[13][4] = 1;	green_platform_transparency_texture[13][5] = 0;	green_platform_transparency_texture[13][6] = 0;	green_platform_transparency_texture[13][7] = 0;	green_platform_transparency_texture[13][8] = 0;	green_platform_transparency_texture[13][9] = 0;	green_platform_transparency_texture[13][10] = 0;	green_platform_transparency_texture[13][11] = 0;	green_platform_transparency_texture[13][12] = 0;	green_platform_transparency_texture[13][13] = 0;	green_platform_transparency_texture[13][14] = 0;	green_platform_transparency_texture[13][15] = 0;	green_platform_transparency_texture[13][16] = 0;	green_platform_transparency_texture[13][17] = 0;	green_platform_transparency_texture[13][18] = 0;	green_platform_transparency_texture[13][19] = 0;	green_platform_transparency_texture[13][20] = 0;	green_platform_transparency_texture[13][21] = 0;	green_platform_transparency_texture[13][22] = 0;	green_platform_transparency_texture[13][23] = 0;	green_platform_transparency_texture[13][24] = 0;	green_platform_transparency_texture[13][25] = 0;	green_platform_transparency_texture[13][26] = 0;	green_platform_transparency_texture[13][27] = 0;	green_platform_transparency_texture[13][28] = 0;	green_platform_transparency_texture[13][29] = 0;	green_platform_transparency_texture[13][30] = 0;	green_platform_transparency_texture[13][31] = 0;	green_platform_transparency_texture[13][32] = 0;	green_platform_transparency_texture[13][33] = 0;	green_platform_transparency_texture[13][34] = 0;	green_platform_transparency_texture[13][35] = 0;	green_platform_transparency_texture[13][36] = 0;	green_platform_transparency_texture[13][37] = 0;	green_platform_transparency_texture[13][38] = 0;	green_platform_transparency_texture[13][39] = 0;	green_platform_transparency_texture[13][40] = 0;	green_platform_transparency_texture[13][41] = 0;	green_platform_transparency_texture[13][42] = 0;	green_platform_transparency_texture[13][43] = 0;	green_platform_transparency_texture[13][44] = 0;	green_platform_transparency_texture[13][45] = 0;	green_platform_transparency_texture[13][46] = 0;	green_platform_transparency_texture[13][47] = 0;	green_platform_transparency_texture[13][48] = 0;	green_platform_transparency_texture[13][49] = 0;	green_platform_transparency_texture[13][50] = 0;	green_platform_transparency_texture[13][51] = 0;	green_platform_transparency_texture[13][52] = 0;	green_platform_transparency_texture[13][53] = 0;	green_platform_transparency_texture[13][54] = 0;	green_platform_transparency_texture[13][55] = 0;	green_platform_transparency_texture[13][56] = 0;	green_platform_transparency_texture[13][57] = 0;	green_platform_transparency_texture[13][58] = 0;	green_platform_transparency_texture[13][59] = 0;	green_platform_transparency_texture[13][60] = 0;	green_platform_transparency_texture[13][61] = 0;	green_platform_transparency_texture[13][62] = 0;	green_platform_transparency_texture[13][63] = 0;	green_platform_transparency_texture[13][64] = 0;	green_platform_transparency_texture[13][65] = 0;	green_platform_transparency_texture[13][66] = 0;	green_platform_transparency_texture[13][67] = 0;	green_platform_transparency_texture[13][68] = 0;	green_platform_transparency_texture[13][69] = 0;	green_platform_transparency_texture[13][70] = 0;	green_platform_transparency_texture[13][71] = 0;	green_platform_transparency_texture[13][72] = 0;	green_platform_transparency_texture[13][73] = 0;	green_platform_transparency_texture[13][74] = 0;	green_platform_transparency_texture[13][75] = 0;	green_platform_transparency_texture[13][76] = 0;	green_platform_transparency_texture[13][77] = 0;	green_platform_transparency_texture[13][78] = 0;	green_platform_transparency_texture[13][79] = 0;	green_platform_transparency_texture[13][80] = 0;	green_platform_transparency_texture[13][81] = 0;	green_platform_transparency_texture[13][82] = 0;	green_platform_transparency_texture[13][83] = 0;	green_platform_transparency_texture[13][84] = 0;	green_platform_transparency_texture[13][85] = 0;	green_platform_transparency_texture[13][86] = 0;	green_platform_transparency_texture[13][87] = 0;	green_platform_transparency_texture[13][88] = 0;	green_platform_transparency_texture[13][89] = 0;	green_platform_transparency_texture[13][90] = 0;	green_platform_transparency_texture[13][91] = 0;	green_platform_transparency_texture[13][92] = 0;	green_platform_transparency_texture[13][93] = 0;	green_platform_transparency_texture[13][94] = 0;	green_platform_transparency_texture[13][95] = 1;	green_platform_transparency_texture[13][96] = 1;	green_platform_transparency_texture[13][97] = 1;	green_platform_transparency_texture[13][98] = 1;	green_platform_transparency_texture[13][99] = 1;	green_platform_transparency_texture[14][0] = 1;	green_platform_transparency_texture[14][1] = 1;	green_platform_transparency_texture[14][2] = 1;	green_platform_transparency_texture[14][3] = 1;	green_platform_transparency_texture[14][4] = 1;	green_platform_transparency_texture[14][5] = 0;	green_platform_transparency_texture[14][6] = 0;	green_platform_transparency_texture[14][7] = 0;	green_platform_transparency_texture[14][8] = 0;	green_platform_transparency_texture[14][9] = 0;	green_platform_transparency_texture[14][10] = 0;	green_platform_transparency_texture[14][11] = 0;	green_platform_transparency_texture[14][12] = 0;	green_platform_transparency_texture[14][13] = 0;	green_platform_transparency_texture[14][14] = 0;	green_platform_transparency_texture[14][15] = 0;	green_platform_transparency_texture[14][16] = 0;	green_platform_transparency_texture[14][17] = 0;	green_platform_transparency_texture[14][18] = 0;	green_platform_transparency_texture[14][19] = 0;	green_platform_transparency_texture[14][20] = 0;	green_platform_transparency_texture[14][21] = 0;	green_platform_transparency_texture[14][22] = 0;	green_platform_transparency_texture[14][23] = 0;	green_platform_transparency_texture[14][24] = 0;	green_platform_transparency_texture[14][25] = 0;	green_platform_transparency_texture[14][26] = 0;	green_platform_transparency_texture[14][27] = 0;	green_platform_transparency_texture[14][28] = 0;	green_platform_transparency_texture[14][29] = 0;	green_platform_transparency_texture[14][30] = 0;	green_platform_transparency_texture[14][31] = 0;	green_platform_transparency_texture[14][32] = 0;	green_platform_transparency_texture[14][33] = 0;	green_platform_transparency_texture[14][34] = 0;	green_platform_transparency_texture[14][35] = 0;	green_platform_transparency_texture[14][36] = 0;	green_platform_transparency_texture[14][37] = 0;	green_platform_transparency_texture[14][38] = 0;	green_platform_transparency_texture[14][39] = 0;	green_platform_transparency_texture[14][40] = 0;	green_platform_transparency_texture[14][41] = 0;	green_platform_transparency_texture[14][42] = 0;	green_platform_transparency_texture[14][43] = 0;	green_platform_transparency_texture[14][44] = 0;	green_platform_transparency_texture[14][45] = 0;	green_platform_transparency_texture[14][46] = 0;	green_platform_transparency_texture[14][47] = 0;	green_platform_transparency_texture[14][48] = 0;	green_platform_transparency_texture[14][49] = 0;	green_platform_transparency_texture[14][50] = 0;	green_platform_transparency_texture[14][51] = 0;	green_platform_transparency_texture[14][52] = 0;	green_platform_transparency_texture[14][53] = 0;	green_platform_transparency_texture[14][54] = 0;	green_platform_transparency_texture[14][55] = 0;	green_platform_transparency_texture[14][56] = 0;	green_platform_transparency_texture[14][57] = 0;	green_platform_transparency_texture[14][58] = 0;	green_platform_transparency_texture[14][59] = 0;	green_platform_transparency_texture[14][60] = 0;	green_platform_transparency_texture[14][61] = 0;	green_platform_transparency_texture[14][62] = 0;	green_platform_transparency_texture[14][63] = 0;	green_platform_transparency_texture[14][64] = 0;	green_platform_transparency_texture[14][65] = 0;	green_platform_transparency_texture[14][66] = 0;	green_platform_transparency_texture[14][67] = 0;	green_platform_transparency_texture[14][68] = 0;	green_platform_transparency_texture[14][69] = 0;	green_platform_transparency_texture[14][70] = 0;	green_platform_transparency_texture[14][71] = 0;	green_platform_transparency_texture[14][72] = 0;	green_platform_transparency_texture[14][73] = 0;	green_platform_transparency_texture[14][74] = 0;	green_platform_transparency_texture[14][75] = 0;	green_platform_transparency_texture[14][76] = 0;	green_platform_transparency_texture[14][77] = 0;	green_platform_transparency_texture[14][78] = 0;	green_platform_transparency_texture[14][79] = 0;	green_platform_transparency_texture[14][80] = 0;	green_platform_transparency_texture[14][81] = 0;	green_platform_transparency_texture[14][82] = 0;	green_platform_transparency_texture[14][83] = 0;	green_platform_transparency_texture[14][84] = 0;	green_platform_transparency_texture[14][85] = 0;	green_platform_transparency_texture[14][86] = 0;	green_platform_transparency_texture[14][87] = 0;	green_platform_transparency_texture[14][88] = 0;	green_platform_transparency_texture[14][89] = 0;	green_platform_transparency_texture[14][90] = 0;	green_platform_transparency_texture[14][91] = 0;	green_platform_transparency_texture[14][92] = 0;	green_platform_transparency_texture[14][93] = 0;	green_platform_transparency_texture[14][94] = 0;	green_platform_transparency_texture[14][95] = 1;	green_platform_transparency_texture[14][96] = 1;	green_platform_transparency_texture[14][97] = 1;	green_platform_transparency_texture[14][98] = 1;	green_platform_transparency_texture[14][99] = 1;	green_platform_transparency_texture[15][0] = 1;	green_platform_transparency_texture[15][1] = 1;	green_platform_transparency_texture[15][2] = 1;	green_platform_transparency_texture[15][3] = 1;	green_platform_transparency_texture[15][4] = 1;	green_platform_transparency_texture[15][5] = 0;	green_platform_transparency_texture[15][6] = 0;	green_platform_transparency_texture[15][7] = 0;	green_platform_transparency_texture[15][8] = 0;	green_platform_transparency_texture[15][9] = 0;	green_platform_transparency_texture[15][10] = 0;	green_platform_transparency_texture[15][11] = 0;	green_platform_transparency_texture[15][12] = 0;	green_platform_transparency_texture[15][13] = 0;	green_platform_transparency_texture[15][14] = 0;	green_platform_transparency_texture[15][15] = 0;	green_platform_transparency_texture[15][16] = 0;	green_platform_transparency_texture[15][17] = 0;	green_platform_transparency_texture[15][18] = 0;	green_platform_transparency_texture[15][19] = 0;	green_platform_transparency_texture[15][20] = 0;	green_platform_transparency_texture[15][21] = 0;	green_platform_transparency_texture[15][22] = 0;	green_platform_transparency_texture[15][23] = 0;	green_platform_transparency_texture[15][24] = 0;	green_platform_transparency_texture[15][25] = 0;	green_platform_transparency_texture[15][26] = 0;	green_platform_transparency_texture[15][27] = 0;	green_platform_transparency_texture[15][28] = 0;	green_platform_transparency_texture[15][29] = 0;	green_platform_transparency_texture[15][30] = 0;	green_platform_transparency_texture[15][31] = 0;	green_platform_transparency_texture[15][32] = 0;	green_platform_transparency_texture[15][33] = 0;	green_platform_transparency_texture[15][34] = 0;	green_platform_transparency_texture[15][35] = 0;	green_platform_transparency_texture[15][36] = 0;	green_platform_transparency_texture[15][37] = 0;	green_platform_transparency_texture[15][38] = 0;	green_platform_transparency_texture[15][39] = 0;	green_platform_transparency_texture[15][40] = 0;	green_platform_transparency_texture[15][41] = 0;	green_platform_transparency_texture[15][42] = 0;	green_platform_transparency_texture[15][43] = 0;	green_platform_transparency_texture[15][44] = 0;	green_platform_transparency_texture[15][45] = 0;	green_platform_transparency_texture[15][46] = 0;	green_platform_transparency_texture[15][47] = 0;	green_platform_transparency_texture[15][48] = 0;	green_platform_transparency_texture[15][49] = 0;	green_platform_transparency_texture[15][50] = 0;	green_platform_transparency_texture[15][51] = 0;	green_platform_transparency_texture[15][52] = 0;	green_platform_transparency_texture[15][53] = 0;	green_platform_transparency_texture[15][54] = 0;	green_platform_transparency_texture[15][55] = 0;	green_platform_transparency_texture[15][56] = 0;	green_platform_transparency_texture[15][57] = 0;	green_platform_transparency_texture[15][58] = 0;	green_platform_transparency_texture[15][59] = 0;	green_platform_transparency_texture[15][60] = 0;	green_platform_transparency_texture[15][61] = 0;	green_platform_transparency_texture[15][62] = 0;	green_platform_transparency_texture[15][63] = 0;	green_platform_transparency_texture[15][64] = 0;	green_platform_transparency_texture[15][65] = 0;	green_platform_transparency_texture[15][66] = 0;	green_platform_transparency_texture[15][67] = 0;	green_platform_transparency_texture[15][68] = 0;	green_platform_transparency_texture[15][69] = 0;	green_platform_transparency_texture[15][70] = 0;	green_platform_transparency_texture[15][71] = 0;	green_platform_transparency_texture[15][72] = 0;	green_platform_transparency_texture[15][73] = 0;	green_platform_transparency_texture[15][74] = 0;	green_platform_transparency_texture[15][75] = 0;	green_platform_transparency_texture[15][76] = 0;	green_platform_transparency_texture[15][77] = 0;	green_platform_transparency_texture[15][78] = 0;	green_platform_transparency_texture[15][79] = 0;	green_platform_transparency_texture[15][80] = 0;	green_platform_transparency_texture[15][81] = 0;	green_platform_transparency_texture[15][82] = 0;	green_platform_transparency_texture[15][83] = 0;	green_platform_transparency_texture[15][84] = 0;	green_platform_transparency_texture[15][85] = 0;	green_platform_transparency_texture[15][86] = 0;	green_platform_transparency_texture[15][87] = 0;	green_platform_transparency_texture[15][88] = 0;	green_platform_transparency_texture[15][89] = 0;	green_platform_transparency_texture[15][90] = 0;	green_platform_transparency_texture[15][91] = 0;	green_platform_transparency_texture[15][92] = 0;	green_platform_transparency_texture[15][93] = 0;	green_platform_transparency_texture[15][94] = 0;	green_platform_transparency_texture[15][95] = 1;	green_platform_transparency_texture[15][96] = 1;	green_platform_transparency_texture[15][97] = 1;	green_platform_transparency_texture[15][98] = 1;	green_platform_transparency_texture[15][99] = 1;	green_platform_transparency_texture[16][0] = 1;	green_platform_transparency_texture[16][1] = 1;	green_platform_transparency_texture[16][2] = 1;	green_platform_transparency_texture[16][3] = 1;	green_platform_transparency_texture[16][4] = 1;	green_platform_transparency_texture[16][5] = 0;	green_platform_transparency_texture[16][6] = 0;	green_platform_transparency_texture[16][7] = 0;	green_platform_transparency_texture[16][8] = 0;	green_platform_transparency_texture[16][9] = 0;	green_platform_transparency_texture[16][10] = 0;	green_platform_transparency_texture[16][11] = 0;	green_platform_transparency_texture[16][12] = 0;	green_platform_transparency_texture[16][13] = 0;	green_platform_transparency_texture[16][14] = 0;	green_platform_transparency_texture[16][15] = 0;	green_platform_transparency_texture[16][16] = 0;	green_platform_transparency_texture[16][17] = 0;	green_platform_transparency_texture[16][18] = 0;	green_platform_transparency_texture[16][19] = 0;	green_platform_transparency_texture[16][20] = 0;	green_platform_transparency_texture[16][21] = 0;	green_platform_transparency_texture[16][22] = 0;	green_platform_transparency_texture[16][23] = 0;	green_platform_transparency_texture[16][24] = 0;	green_platform_transparency_texture[16][25] = 0;	green_platform_transparency_texture[16][26] = 0;	green_platform_transparency_texture[16][27] = 0;	green_platform_transparency_texture[16][28] = 0;	green_platform_transparency_texture[16][29] = 0;	green_platform_transparency_texture[16][30] = 0;	green_platform_transparency_texture[16][31] = 0;	green_platform_transparency_texture[16][32] = 0;	green_platform_transparency_texture[16][33] = 0;	green_platform_transparency_texture[16][34] = 0;	green_platform_transparency_texture[16][35] = 0;	green_platform_transparency_texture[16][36] = 0;	green_platform_transparency_texture[16][37] = 0;	green_platform_transparency_texture[16][38] = 0;	green_platform_transparency_texture[16][39] = 0;	green_platform_transparency_texture[16][40] = 0;	green_platform_transparency_texture[16][41] = 0;	green_platform_transparency_texture[16][42] = 0;	green_platform_transparency_texture[16][43] = 0;	green_platform_transparency_texture[16][44] = 0;	green_platform_transparency_texture[16][45] = 0;	green_platform_transparency_texture[16][46] = 0;	green_platform_transparency_texture[16][47] = 0;	green_platform_transparency_texture[16][48] = 0;	green_platform_transparency_texture[16][49] = 0;	green_platform_transparency_texture[16][50] = 0;	green_platform_transparency_texture[16][51] = 0;	green_platform_transparency_texture[16][52] = 0;	green_platform_transparency_texture[16][53] = 0;	green_platform_transparency_texture[16][54] = 0;	green_platform_transparency_texture[16][55] = 0;	green_platform_transparency_texture[16][56] = 0;	green_platform_transparency_texture[16][57] = 0;	green_platform_transparency_texture[16][58] = 0;	green_platform_transparency_texture[16][59] = 0;	green_platform_transparency_texture[16][60] = 0;	green_platform_transparency_texture[16][61] = 0;	green_platform_transparency_texture[16][62] = 0;	green_platform_transparency_texture[16][63] = 0;	green_platform_transparency_texture[16][64] = 0;	green_platform_transparency_texture[16][65] = 0;	green_platform_transparency_texture[16][66] = 0;	green_platform_transparency_texture[16][67] = 0;	green_platform_transparency_texture[16][68] = 0;	green_platform_transparency_texture[16][69] = 0;	green_platform_transparency_texture[16][70] = 0;	green_platform_transparency_texture[16][71] = 0;	green_platform_transparency_texture[16][72] = 0;	green_platform_transparency_texture[16][73] = 0;	green_platform_transparency_texture[16][74] = 0;	green_platform_transparency_texture[16][75] = 0;	green_platform_transparency_texture[16][76] = 0;	green_platform_transparency_texture[16][77] = 0;	green_platform_transparency_texture[16][78] = 0;	green_platform_transparency_texture[16][79] = 0;	green_platform_transparency_texture[16][80] = 0;	green_platform_transparency_texture[16][81] = 0;	green_platform_transparency_texture[16][82] = 0;	green_platform_transparency_texture[16][83] = 0;	green_platform_transparency_texture[16][84] = 0;	green_platform_transparency_texture[16][85] = 0;	green_platform_transparency_texture[16][86] = 0;	green_platform_transparency_texture[16][87] = 0;	green_platform_transparency_texture[16][88] = 0;	green_platform_transparency_texture[16][89] = 0;	green_platform_transparency_texture[16][90] = 0;	green_platform_transparency_texture[16][91] = 0;	green_platform_transparency_texture[16][92] = 0;	green_platform_transparency_texture[16][93] = 0;	green_platform_transparency_texture[16][94] = 0;	green_platform_transparency_texture[16][95] = 1;	green_platform_transparency_texture[16][96] = 1;	green_platform_transparency_texture[16][97] = 1;	green_platform_transparency_texture[16][98] = 1;	green_platform_transparency_texture[16][99] = 1;	green_platform_transparency_texture[17][0] = 1;	green_platform_transparency_texture[17][1] = 1;	green_platform_transparency_texture[17][2] = 1;	green_platform_transparency_texture[17][3] = 1;	green_platform_transparency_texture[17][4] = 1;	green_platform_transparency_texture[17][5] = 0;	green_platform_transparency_texture[17][6] = 0;	green_platform_transparency_texture[17][7] = 0;	green_platform_transparency_texture[17][8] = 0;	green_platform_transparency_texture[17][9] = 0;	green_platform_transparency_texture[17][10] = 0;	green_platform_transparency_texture[17][11] = 0;	green_platform_transparency_texture[17][12] = 0;	green_platform_transparency_texture[17][13] = 0;	green_platform_transparency_texture[17][14] = 0;	green_platform_transparency_texture[17][15] = 0;	green_platform_transparency_texture[17][16] = 0;	green_platform_transparency_texture[17][17] = 0;	green_platform_transparency_texture[17][18] = 0;	green_platform_transparency_texture[17][19] = 0;	green_platform_transparency_texture[17][20] = 0;	green_platform_transparency_texture[17][21] = 0;	green_platform_transparency_texture[17][22] = 0;	green_platform_transparency_texture[17][23] = 0;	green_platform_transparency_texture[17][24] = 0;	green_platform_transparency_texture[17][25] = 0;	green_platform_transparency_texture[17][26] = 0;	green_platform_transparency_texture[17][27] = 0;	green_platform_transparency_texture[17][28] = 0;	green_platform_transparency_texture[17][29] = 0;	green_platform_transparency_texture[17][30] = 0;	green_platform_transparency_texture[17][31] = 0;	green_platform_transparency_texture[17][32] = 0;	green_platform_transparency_texture[17][33] = 0;	green_platform_transparency_texture[17][34] = 0;	green_platform_transparency_texture[17][35] = 0;	green_platform_transparency_texture[17][36] = 0;	green_platform_transparency_texture[17][37] = 0;	green_platform_transparency_texture[17][38] = 0;	green_platform_transparency_texture[17][39] = 0;	green_platform_transparency_texture[17][40] = 0;	green_platform_transparency_texture[17][41] = 0;	green_platform_transparency_texture[17][42] = 0;	green_platform_transparency_texture[17][43] = 0;	green_platform_transparency_texture[17][44] = 0;	green_platform_transparency_texture[17][45] = 0;	green_platform_transparency_texture[17][46] = 0;	green_platform_transparency_texture[17][47] = 0;	green_platform_transparency_texture[17][48] = 0;	green_platform_transparency_texture[17][49] = 0;	green_platform_transparency_texture[17][50] = 0;	green_platform_transparency_texture[17][51] = 0;	green_platform_transparency_texture[17][52] = 0;	green_platform_transparency_texture[17][53] = 0;	green_platform_transparency_texture[17][54] = 0;	green_platform_transparency_texture[17][55] = 0;	green_platform_transparency_texture[17][56] = 0;	green_platform_transparency_texture[17][57] = 0;	green_platform_transparency_texture[17][58] = 0;	green_platform_transparency_texture[17][59] = 0;	green_platform_transparency_texture[17][60] = 0;	green_platform_transparency_texture[17][61] = 0;	green_platform_transparency_texture[17][62] = 0;	green_platform_transparency_texture[17][63] = 0;	green_platform_transparency_texture[17][64] = 0;	green_platform_transparency_texture[17][65] = 0;	green_platform_transparency_texture[17][66] = 0;	green_platform_transparency_texture[17][67] = 0;	green_platform_transparency_texture[17][68] = 0;	green_platform_transparency_texture[17][69] = 0;	green_platform_transparency_texture[17][70] = 0;	green_platform_transparency_texture[17][71] = 0;	green_platform_transparency_texture[17][72] = 0;	green_platform_transparency_texture[17][73] = 0;	green_platform_transparency_texture[17][74] = 0;	green_platform_transparency_texture[17][75] = 0;	green_platform_transparency_texture[17][76] = 0;	green_platform_transparency_texture[17][77] = 0;	green_platform_transparency_texture[17][78] = 0;	green_platform_transparency_texture[17][79] = 0;	green_platform_transparency_texture[17][80] = 0;	green_platform_transparency_texture[17][81] = 0;	green_platform_transparency_texture[17][82] = 0;	green_platform_transparency_texture[17][83] = 0;	green_platform_transparency_texture[17][84] = 0;	green_platform_transparency_texture[17][85] = 0;	green_platform_transparency_texture[17][86] = 0;	green_platform_transparency_texture[17][87] = 0;	green_platform_transparency_texture[17][88] = 0;	green_platform_transparency_texture[17][89] = 0;	green_platform_transparency_texture[17][90] = 0;	green_platform_transparency_texture[17][91] = 0;	green_platform_transparency_texture[17][92] = 0;	green_platform_transparency_texture[17][93] = 0;	green_platform_transparency_texture[17][94] = 0;	green_platform_transparency_texture[17][95] = 1;	green_platform_transparency_texture[17][96] = 1;	green_platform_transparency_texture[17][97] = 1;	green_platform_transparency_texture[17][98] = 1;	green_platform_transparency_texture[17][99] = 1;	green_platform_transparency_texture[18][0] = 1;	green_platform_transparency_texture[18][1] = 1;	green_platform_transparency_texture[18][2] = 1;	green_platform_transparency_texture[18][3] = 1;	green_platform_transparency_texture[18][4] = 1;	green_platform_transparency_texture[18][5] = 0;	green_platform_transparency_texture[18][6] = 0;	green_platform_transparency_texture[18][7] = 0;	green_platform_transparency_texture[18][8] = 0;	green_platform_transparency_texture[18][9] = 0;	green_platform_transparency_texture[18][10] = 0;	green_platform_transparency_texture[18][11] = 0;	green_platform_transparency_texture[18][12] = 0;	green_platform_transparency_texture[18][13] = 0;	green_platform_transparency_texture[18][14] = 0;	green_platform_transparency_texture[18][15] = 0;	green_platform_transparency_texture[18][16] = 0;	green_platform_transparency_texture[18][17] = 0;	green_platform_transparency_texture[18][18] = 0;	green_platform_transparency_texture[18][19] = 0;	green_platform_transparency_texture[18][20] = 0;	green_platform_transparency_texture[18][21] = 0;	green_platform_transparency_texture[18][22] = 0;	green_platform_transparency_texture[18][23] = 0;	green_platform_transparency_texture[18][24] = 0;	green_platform_transparency_texture[18][25] = 0;	green_platform_transparency_texture[18][26] = 0;	green_platform_transparency_texture[18][27] = 0;	green_platform_transparency_texture[18][28] = 0;	green_platform_transparency_texture[18][29] = 0;	green_platform_transparency_texture[18][30] = 0;	green_platform_transparency_texture[18][31] = 0;	green_platform_transparency_texture[18][32] = 0;	green_platform_transparency_texture[18][33] = 0;	green_platform_transparency_texture[18][34] = 0;	green_platform_transparency_texture[18][35] = 0;	green_platform_transparency_texture[18][36] = 0;	green_platform_transparency_texture[18][37] = 0;	green_platform_transparency_texture[18][38] = 0;	green_platform_transparency_texture[18][39] = 0;	green_platform_transparency_texture[18][40] = 0;	green_platform_transparency_texture[18][41] = 0;	green_platform_transparency_texture[18][42] = 0;	green_platform_transparency_texture[18][43] = 0;	green_platform_transparency_texture[18][44] = 0;	green_platform_transparency_texture[18][45] = 0;	green_platform_transparency_texture[18][46] = 0;	green_platform_transparency_texture[18][47] = 0;	green_platform_transparency_texture[18][48] = 0;	green_platform_transparency_texture[18][49] = 0;	green_platform_transparency_texture[18][50] = 0;	green_platform_transparency_texture[18][51] = 0;	green_platform_transparency_texture[18][52] = 0;	green_platform_transparency_texture[18][53] = 0;	green_platform_transparency_texture[18][54] = 0;	green_platform_transparency_texture[18][55] = 0;	green_platform_transparency_texture[18][56] = 0;	green_platform_transparency_texture[18][57] = 0;	green_platform_transparency_texture[18][58] = 0;	green_platform_transparency_texture[18][59] = 0;	green_platform_transparency_texture[18][60] = 0;	green_platform_transparency_texture[18][61] = 0;	green_platform_transparency_texture[18][62] = 0;	green_platform_transparency_texture[18][63] = 0;	green_platform_transparency_texture[18][64] = 0;	green_platform_transparency_texture[18][65] = 0;	green_platform_transparency_texture[18][66] = 0;	green_platform_transparency_texture[18][67] = 0;	green_platform_transparency_texture[18][68] = 0;	green_platform_transparency_texture[18][69] = 0;	green_platform_transparency_texture[18][70] = 0;	green_platform_transparency_texture[18][71] = 0;	green_platform_transparency_texture[18][72] = 0;	green_platform_transparency_texture[18][73] = 0;	green_platform_transparency_texture[18][74] = 0;	green_platform_transparency_texture[18][75] = 0;	green_platform_transparency_texture[18][76] = 0;	green_platform_transparency_texture[18][77] = 0;	green_platform_transparency_texture[18][78] = 0;	green_platform_transparency_texture[18][79] = 0;	green_platform_transparency_texture[18][80] = 0;	green_platform_transparency_texture[18][81] = 0;	green_platform_transparency_texture[18][82] = 0;	green_platform_transparency_texture[18][83] = 0;	green_platform_transparency_texture[18][84] = 0;	green_platform_transparency_texture[18][85] = 0;	green_platform_transparency_texture[18][86] = 0;	green_platform_transparency_texture[18][87] = 0;	green_platform_transparency_texture[18][88] = 0;	green_platform_transparency_texture[18][89] = 0;	green_platform_transparency_texture[18][90] = 0;	green_platform_transparency_texture[18][91] = 0;	green_platform_transparency_texture[18][92] = 0;	green_platform_transparency_texture[18][93] = 0;	green_platform_transparency_texture[18][94] = 0;	green_platform_transparency_texture[18][95] = 1;	green_platform_transparency_texture[18][96] = 1;	green_platform_transparency_texture[18][97] = 1;	green_platform_transparency_texture[18][98] = 1;	green_platform_transparency_texture[18][99] = 1;	green_platform_transparency_texture[19][0] = 1;	green_platform_transparency_texture[19][1] = 1;	green_platform_transparency_texture[19][2] = 1;	green_platform_transparency_texture[19][3] = 1;	green_platform_transparency_texture[19][4] = 1;	green_platform_transparency_texture[19][5] = 0;	green_platform_transparency_texture[19][6] = 0;	green_platform_transparency_texture[19][7] = 0;	green_platform_transparency_texture[19][8] = 0;	green_platform_transparency_texture[19][9] = 0;	green_platform_transparency_texture[19][10] = 0;	green_platform_transparency_texture[19][11] = 0;	green_platform_transparency_texture[19][12] = 0;	green_platform_transparency_texture[19][13] = 0;	green_platform_transparency_texture[19][14] = 0;	green_platform_transparency_texture[19][15] = 0;	green_platform_transparency_texture[19][16] = 0;	green_platform_transparency_texture[19][17] = 0;	green_platform_transparency_texture[19][18] = 0;	green_platform_transparency_texture[19][19] = 0;	green_platform_transparency_texture[19][20] = 0;	green_platform_transparency_texture[19][21] = 0;	green_platform_transparency_texture[19][22] = 0;	green_platform_transparency_texture[19][23] = 0;	green_platform_transparency_texture[19][24] = 0;	green_platform_transparency_texture[19][25] = 0;	green_platform_transparency_texture[19][26] = 0;	green_platform_transparency_texture[19][27] = 0;	green_platform_transparency_texture[19][28] = 0;	green_platform_transparency_texture[19][29] = 0;	green_platform_transparency_texture[19][30] = 0;	green_platform_transparency_texture[19][31] = 0;	green_platform_transparency_texture[19][32] = 0;	green_platform_transparency_texture[19][33] = 0;	green_platform_transparency_texture[19][34] = 0;	green_platform_transparency_texture[19][35] = 0;	green_platform_transparency_texture[19][36] = 0;	green_platform_transparency_texture[19][37] = 0;	green_platform_transparency_texture[19][38] = 0;	green_platform_transparency_texture[19][39] = 0;	green_platform_transparency_texture[19][40] = 0;	green_platform_transparency_texture[19][41] = 0;	green_platform_transparency_texture[19][42] = 0;	green_platform_transparency_texture[19][43] = 0;	green_platform_transparency_texture[19][44] = 0;	green_platform_transparency_texture[19][45] = 0;	green_platform_transparency_texture[19][46] = 0;	green_platform_transparency_texture[19][47] = 0;	green_platform_transparency_texture[19][48] = 0;	green_platform_transparency_texture[19][49] = 0;	green_platform_transparency_texture[19][50] = 0;	green_platform_transparency_texture[19][51] = 0;	green_platform_transparency_texture[19][52] = 0;	green_platform_transparency_texture[19][53] = 0;	green_platform_transparency_texture[19][54] = 0;	green_platform_transparency_texture[19][55] = 0;	green_platform_transparency_texture[19][56] = 0;	green_platform_transparency_texture[19][57] = 0;	green_platform_transparency_texture[19][58] = 0;	green_platform_transparency_texture[19][59] = 0;	green_platform_transparency_texture[19][60] = 0;	green_platform_transparency_texture[19][61] = 0;	green_platform_transparency_texture[19][62] = 0;	green_platform_transparency_texture[19][63] = 0;	green_platform_transparency_texture[19][64] = 0;	green_platform_transparency_texture[19][65] = 0;	green_platform_transparency_texture[19][66] = 0;	green_platform_transparency_texture[19][67] = 0;	green_platform_transparency_texture[19][68] = 0;	green_platform_transparency_texture[19][69] = 0;	green_platform_transparency_texture[19][70] = 0;	green_platform_transparency_texture[19][71] = 0;	green_platform_transparency_texture[19][72] = 0;	green_platform_transparency_texture[19][73] = 0;	green_platform_transparency_texture[19][74] = 0;	green_platform_transparency_texture[19][75] = 0;	green_platform_transparency_texture[19][76] = 0;	green_platform_transparency_texture[19][77] = 0;	green_platform_transparency_texture[19][78] = 0;	green_platform_transparency_texture[19][79] = 0;	green_platform_transparency_texture[19][80] = 0;	green_platform_transparency_texture[19][81] = 0;	green_platform_transparency_texture[19][82] = 0;	green_platform_transparency_texture[19][83] = 0;	green_platform_transparency_texture[19][84] = 0;	green_platform_transparency_texture[19][85] = 0;	green_platform_transparency_texture[19][86] = 0;	green_platform_transparency_texture[19][87] = 0;	green_platform_transparency_texture[19][88] = 0;	green_platform_transparency_texture[19][89] = 0;	green_platform_transparency_texture[19][90] = 0;	green_platform_transparency_texture[19][91] = 0;	green_platform_transparency_texture[19][92] = 0;	green_platform_transparency_texture[19][93] = 0;	green_platform_transparency_texture[19][94] = 0;	green_platform_transparency_texture[19][95] = 1;	green_platform_transparency_texture[19][96] = 1;	green_platform_transparency_texture[19][97] = 1;	green_platform_transparency_texture[19][98] = 1;	green_platform_transparency_texture[19][99] = 1;	green_platform_transparency_texture[20][0] = 1;	green_platform_transparency_texture[20][1] = 1;	green_platform_transparency_texture[20][2] = 1;	green_platform_transparency_texture[20][3] = 1;	green_platform_transparency_texture[20][4] = 1;	green_platform_transparency_texture[20][5] = 1;	green_platform_transparency_texture[20][6] = 1;	green_platform_transparency_texture[20][7] = 1;	green_platform_transparency_texture[20][8] = 1;	green_platform_transparency_texture[20][9] = 0;	green_platform_transparency_texture[20][10] = 0;	green_platform_transparency_texture[20][11] = 0;	green_platform_transparency_texture[20][12] = 0;	green_platform_transparency_texture[20][13] = 0;	green_platform_transparency_texture[20][14] = 0;	green_platform_transparency_texture[20][15] = 0;	green_platform_transparency_texture[20][16] = 0;	green_platform_transparency_texture[20][17] = 0;	green_platform_transparency_texture[20][18] = 0;	green_platform_transparency_texture[20][19] = 0;	green_platform_transparency_texture[20][20] = 0;	green_platform_transparency_texture[20][21] = 0;	green_platform_transparency_texture[20][22] = 0;	green_platform_transparency_texture[20][23] = 0;	green_platform_transparency_texture[20][24] = 0;	green_platform_transparency_texture[20][25] = 0;	green_platform_transparency_texture[20][26] = 0;	green_platform_transparency_texture[20][27] = 0;	green_platform_transparency_texture[20][28] = 0;	green_platform_transparency_texture[20][29] = 0;	green_platform_transparency_texture[20][30] = 0;	green_platform_transparency_texture[20][31] = 0;	green_platform_transparency_texture[20][32] = 0;	green_platform_transparency_texture[20][33] = 0;	green_platform_transparency_texture[20][34] = 0;	green_platform_transparency_texture[20][35] = 0;	green_platform_transparency_texture[20][36] = 0;	green_platform_transparency_texture[20][37] = 0;	green_platform_transparency_texture[20][38] = 0;	green_platform_transparency_texture[20][39] = 0;	green_platform_transparency_texture[20][40] = 0;	green_platform_transparency_texture[20][41] = 0;	green_platform_transparency_texture[20][42] = 0;	green_platform_transparency_texture[20][43] = 0;	green_platform_transparency_texture[20][44] = 0;	green_platform_transparency_texture[20][45] = 0;	green_platform_transparency_texture[20][46] = 0;	green_platform_transparency_texture[20][47] = 0;	green_platform_transparency_texture[20][48] = 0;	green_platform_transparency_texture[20][49] = 0;	green_platform_transparency_texture[20][50] = 0;	green_platform_transparency_texture[20][51] = 0;	green_platform_transparency_texture[20][52] = 0;	green_platform_transparency_texture[20][53] = 0;	green_platform_transparency_texture[20][54] = 0;	green_platform_transparency_texture[20][55] = 0;	green_platform_transparency_texture[20][56] = 0;	green_platform_transparency_texture[20][57] = 0;	green_platform_transparency_texture[20][58] = 0;	green_platform_transparency_texture[20][59] = 0;	green_platform_transparency_texture[20][60] = 0;	green_platform_transparency_texture[20][61] = 0;	green_platform_transparency_texture[20][62] = 0;	green_platform_transparency_texture[20][63] = 0;	green_platform_transparency_texture[20][64] = 0;	green_platform_transparency_texture[20][65] = 0;	green_platform_transparency_texture[20][66] = 0;	green_platform_transparency_texture[20][67] = 0;	green_platform_transparency_texture[20][68] = 0;	green_platform_transparency_texture[20][69] = 0;	green_platform_transparency_texture[20][70] = 0;	green_platform_transparency_texture[20][71] = 0;	green_platform_transparency_texture[20][72] = 0;	green_platform_transparency_texture[20][73] = 0;	green_platform_transparency_texture[20][74] = 0;	green_platform_transparency_texture[20][75] = 0;	green_platform_transparency_texture[20][76] = 0;	green_platform_transparency_texture[20][77] = 0;	green_platform_transparency_texture[20][78] = 0;	green_platform_transparency_texture[20][79] = 0;	green_platform_transparency_texture[20][80] = 0;	green_platform_transparency_texture[20][81] = 0;	green_platform_transparency_texture[20][82] = 0;	green_platform_transparency_texture[20][83] = 0;	green_platform_transparency_texture[20][84] = 0;	green_platform_transparency_texture[20][85] = 0;	green_platform_transparency_texture[20][86] = 0;	green_platform_transparency_texture[20][87] = 0;	green_platform_transparency_texture[20][88] = 0;	green_platform_transparency_texture[20][89] = 0;	green_platform_transparency_texture[20][90] = 1;	green_platform_transparency_texture[20][91] = 1;	green_platform_transparency_texture[20][92] = 1;	green_platform_transparency_texture[20][93] = 1;	green_platform_transparency_texture[20][94] = 1;	green_platform_transparency_texture[20][95] = 1;	green_platform_transparency_texture[20][96] = 1;	green_platform_transparency_texture[20][97] = 1;	green_platform_transparency_texture[20][98] = 1;	green_platform_transparency_texture[20][99] = 1;	green_platform_transparency_texture[21][0] = 1;	green_platform_transparency_texture[21][1] = 1;	green_platform_transparency_texture[21][2] = 1;	green_platform_transparency_texture[21][3] = 1;	green_platform_transparency_texture[21][4] = 1;	green_platform_transparency_texture[21][5] = 1;	green_platform_transparency_texture[21][6] = 1;	green_platform_transparency_texture[21][7] = 1;	green_platform_transparency_texture[21][8] = 1;	green_platform_transparency_texture[21][9] = 0;	green_platform_transparency_texture[21][10] = 0;	green_platform_transparency_texture[21][11] = 0;	green_platform_transparency_texture[21][12] = 0;	green_platform_transparency_texture[21][13] = 0;	green_platform_transparency_texture[21][14] = 0;	green_platform_transparency_texture[21][15] = 0;	green_platform_transparency_texture[21][16] = 0;	green_platform_transparency_texture[21][17] = 0;	green_platform_transparency_texture[21][18] = 0;	green_platform_transparency_texture[21][19] = 0;	green_platform_transparency_texture[21][20] = 0;	green_platform_transparency_texture[21][21] = 0;	green_platform_transparency_texture[21][22] = 0;	green_platform_transparency_texture[21][23] = 0;	green_platform_transparency_texture[21][24] = 0;	green_platform_transparency_texture[21][25] = 0;	green_platform_transparency_texture[21][26] = 0;	green_platform_transparency_texture[21][27] = 0;	green_platform_transparency_texture[21][28] = 0;	green_platform_transparency_texture[21][29] = 0;	green_platform_transparency_texture[21][30] = 0;	green_platform_transparency_texture[21][31] = 0;	green_platform_transparency_texture[21][32] = 0;	green_platform_transparency_texture[21][33] = 0;	green_platform_transparency_texture[21][34] = 0;	green_platform_transparency_texture[21][35] = 0;	green_platform_transparency_texture[21][36] = 0;	green_platform_transparency_texture[21][37] = 0;	green_platform_transparency_texture[21][38] = 0;	green_platform_transparency_texture[21][39] = 0;	green_platform_transparency_texture[21][40] = 0;	green_platform_transparency_texture[21][41] = 0;	green_platform_transparency_texture[21][42] = 0;	green_platform_transparency_texture[21][43] = 0;	green_platform_transparency_texture[21][44] = 0;	green_platform_transparency_texture[21][45] = 0;	green_platform_transparency_texture[21][46] = 0;	green_platform_transparency_texture[21][47] = 0;	green_platform_transparency_texture[21][48] = 0;	green_platform_transparency_texture[21][49] = 0;	green_platform_transparency_texture[21][50] = 0;	green_platform_transparency_texture[21][51] = 0;	green_platform_transparency_texture[21][52] = 0;	green_platform_transparency_texture[21][53] = 0;	green_platform_transparency_texture[21][54] = 0;	green_platform_transparency_texture[21][55] = 0;	green_platform_transparency_texture[21][56] = 0;	green_platform_transparency_texture[21][57] = 0;	green_platform_transparency_texture[21][58] = 0;	green_platform_transparency_texture[21][59] = 0;	green_platform_transparency_texture[21][60] = 0;	green_platform_transparency_texture[21][61] = 0;	green_platform_transparency_texture[21][62] = 0;	green_platform_transparency_texture[21][63] = 0;	green_platform_transparency_texture[21][64] = 0;	green_platform_transparency_texture[21][65] = 0;	green_platform_transparency_texture[21][66] = 0;	green_platform_transparency_texture[21][67] = 0;	green_platform_transparency_texture[21][68] = 0;	green_platform_transparency_texture[21][69] = 0;	green_platform_transparency_texture[21][70] = 0;	green_platform_transparency_texture[21][71] = 0;	green_platform_transparency_texture[21][72] = 0;	green_platform_transparency_texture[21][73] = 0;	green_platform_transparency_texture[21][74] = 0;	green_platform_transparency_texture[21][75] = 0;	green_platform_transparency_texture[21][76] = 0;	green_platform_transparency_texture[21][77] = 0;	green_platform_transparency_texture[21][78] = 0;	green_platform_transparency_texture[21][79] = 0;	green_platform_transparency_texture[21][80] = 0;	green_platform_transparency_texture[21][81] = 0;	green_platform_transparency_texture[21][82] = 0;	green_platform_transparency_texture[21][83] = 0;	green_platform_transparency_texture[21][84] = 0;	green_platform_transparency_texture[21][85] = 0;	green_platform_transparency_texture[21][86] = 0;	green_platform_transparency_texture[21][87] = 0;	green_platform_transparency_texture[21][88] = 0;	green_platform_transparency_texture[21][89] = 0;	green_platform_transparency_texture[21][90] = 1;	green_platform_transparency_texture[21][91] = 1;	green_platform_transparency_texture[21][92] = 1;	green_platform_transparency_texture[21][93] = 1;	green_platform_transparency_texture[21][94] = 1;	green_platform_transparency_texture[21][95] = 1;	green_platform_transparency_texture[21][96] = 1;	green_platform_transparency_texture[21][97] = 1;	green_platform_transparency_texture[21][98] = 1;	green_platform_transparency_texture[21][99] = 1;	green_platform_transparency_texture[22][0] = 1;	green_platform_transparency_texture[22][1] = 1;	green_platform_transparency_texture[22][2] = 1;	green_platform_transparency_texture[22][3] = 1;	green_platform_transparency_texture[22][4] = 1;	green_platform_transparency_texture[22][5] = 1;	green_platform_transparency_texture[22][6] = 1;	green_platform_transparency_texture[22][7] = 1;	green_platform_transparency_texture[22][8] = 1;	green_platform_transparency_texture[22][9] = 0;	green_platform_transparency_texture[22][10] = 0;	green_platform_transparency_texture[22][11] = 0;	green_platform_transparency_texture[22][12] = 0;	green_platform_transparency_texture[22][13] = 0;	green_platform_transparency_texture[22][14] = 0;	green_platform_transparency_texture[22][15] = 0;	green_platform_transparency_texture[22][16] = 0;	green_platform_transparency_texture[22][17] = 0;	green_platform_transparency_texture[22][18] = 0;	green_platform_transparency_texture[22][19] = 0;	green_platform_transparency_texture[22][20] = 0;	green_platform_transparency_texture[22][21] = 0;	green_platform_transparency_texture[22][22] = 0;	green_platform_transparency_texture[22][23] = 0;	green_platform_transparency_texture[22][24] = 0;	green_platform_transparency_texture[22][25] = 0;	green_platform_transparency_texture[22][26] = 0;	green_platform_transparency_texture[22][27] = 0;	green_platform_transparency_texture[22][28] = 0;	green_platform_transparency_texture[22][29] = 0;	green_platform_transparency_texture[22][30] = 0;	green_platform_transparency_texture[22][31] = 0;	green_platform_transparency_texture[22][32] = 0;	green_platform_transparency_texture[22][33] = 0;	green_platform_transparency_texture[22][34] = 0;	green_platform_transparency_texture[22][35] = 0;	green_platform_transparency_texture[22][36] = 0;	green_platform_transparency_texture[22][37] = 0;	green_platform_transparency_texture[22][38] = 0;	green_platform_transparency_texture[22][39] = 0;	green_platform_transparency_texture[22][40] = 0;	green_platform_transparency_texture[22][41] = 0;	green_platform_transparency_texture[22][42] = 0;	green_platform_transparency_texture[22][43] = 0;	green_platform_transparency_texture[22][44] = 0;	green_platform_transparency_texture[22][45] = 0;	green_platform_transparency_texture[22][46] = 0;	green_platform_transparency_texture[22][47] = 0;	green_platform_transparency_texture[22][48] = 0;	green_platform_transparency_texture[22][49] = 0;	green_platform_transparency_texture[22][50] = 0;	green_platform_transparency_texture[22][51] = 0;	green_platform_transparency_texture[22][52] = 0;	green_platform_transparency_texture[22][53] = 0;	green_platform_transparency_texture[22][54] = 0;	green_platform_transparency_texture[22][55] = 0;	green_platform_transparency_texture[22][56] = 0;	green_platform_transparency_texture[22][57] = 0;	green_platform_transparency_texture[22][58] = 0;	green_platform_transparency_texture[22][59] = 0;	green_platform_transparency_texture[22][60] = 0;	green_platform_transparency_texture[22][61] = 0;	green_platform_transparency_texture[22][62] = 0;	green_platform_transparency_texture[22][63] = 0;	green_platform_transparency_texture[22][64] = 0;	green_platform_transparency_texture[22][65] = 0;	green_platform_transparency_texture[22][66] = 0;	green_platform_transparency_texture[22][67] = 0;	green_platform_transparency_texture[22][68] = 0;	green_platform_transparency_texture[22][69] = 0;	green_platform_transparency_texture[22][70] = 0;	green_platform_transparency_texture[22][71] = 0;	green_platform_transparency_texture[22][72] = 0;	green_platform_transparency_texture[22][73] = 0;	green_platform_transparency_texture[22][74] = 0;	green_platform_transparency_texture[22][75] = 0;	green_platform_transparency_texture[22][76] = 0;	green_platform_transparency_texture[22][77] = 0;	green_platform_transparency_texture[22][78] = 0;	green_platform_transparency_texture[22][79] = 0;	green_platform_transparency_texture[22][80] = 0;	green_platform_transparency_texture[22][81] = 0;	green_platform_transparency_texture[22][82] = 0;	green_platform_transparency_texture[22][83] = 0;	green_platform_transparency_texture[22][84] = 0;	green_platform_transparency_texture[22][85] = 0;	green_platform_transparency_texture[22][86] = 0;	green_platform_transparency_texture[22][87] = 0;	green_platform_transparency_texture[22][88] = 0;	green_platform_transparency_texture[22][89] = 0;	green_platform_transparency_texture[22][90] = 1;	green_platform_transparency_texture[22][91] = 1;	green_platform_transparency_texture[22][92] = 1;	green_platform_transparency_texture[22][93] = 1;	green_platform_transparency_texture[22][94] = 1;	green_platform_transparency_texture[22][95] = 1;	green_platform_transparency_texture[22][96] = 1;	green_platform_transparency_texture[22][97] = 1;	green_platform_transparency_texture[22][98] = 1;	green_platform_transparency_texture[22][99] = 1;	green_platform_transparency_texture[23][0] = 1;	green_platform_transparency_texture[23][1] = 1;	green_platform_transparency_texture[23][2] = 1;	green_platform_transparency_texture[23][3] = 1;	green_platform_transparency_texture[23][4] = 1;	green_platform_transparency_texture[23][5] = 1;	green_platform_transparency_texture[23][6] = 1;	green_platform_transparency_texture[23][7] = 1;	green_platform_transparency_texture[23][8] = 1;	green_platform_transparency_texture[23][9] = 0;	green_platform_transparency_texture[23][10] = 0;	green_platform_transparency_texture[23][11] = 0;	green_platform_transparency_texture[23][12] = 0;	green_platform_transparency_texture[23][13] = 0;	green_platform_transparency_texture[23][14] = 0;	green_platform_transparency_texture[23][15] = 0;	green_platform_transparency_texture[23][16] = 0;	green_platform_transparency_texture[23][17] = 0;	green_platform_transparency_texture[23][18] = 0;	green_platform_transparency_texture[23][19] = 0;	green_platform_transparency_texture[23][20] = 0;	green_platform_transparency_texture[23][21] = 0;	green_platform_transparency_texture[23][22] = 0;	green_platform_transparency_texture[23][23] = 0;	green_platform_transparency_texture[23][24] = 0;	green_platform_transparency_texture[23][25] = 0;	green_platform_transparency_texture[23][26] = 0;	green_platform_transparency_texture[23][27] = 0;	green_platform_transparency_texture[23][28] = 0;	green_platform_transparency_texture[23][29] = 0;	green_platform_transparency_texture[23][30] = 0;	green_platform_transparency_texture[23][31] = 0;	green_platform_transparency_texture[23][32] = 0;	green_platform_transparency_texture[23][33] = 0;	green_platform_transparency_texture[23][34] = 0;	green_platform_transparency_texture[23][35] = 0;	green_platform_transparency_texture[23][36] = 0;	green_platform_transparency_texture[23][37] = 0;	green_platform_transparency_texture[23][38] = 0;	green_platform_transparency_texture[23][39] = 0;	green_platform_transparency_texture[23][40] = 0;	green_platform_transparency_texture[23][41] = 0;	green_platform_transparency_texture[23][42] = 0;	green_platform_transparency_texture[23][43] = 0;	green_platform_transparency_texture[23][44] = 0;	green_platform_transparency_texture[23][45] = 0;	green_platform_transparency_texture[23][46] = 0;	green_platform_transparency_texture[23][47] = 0;	green_platform_transparency_texture[23][48] = 0;	green_platform_transparency_texture[23][49] = 0;	green_platform_transparency_texture[23][50] = 0;	green_platform_transparency_texture[23][51] = 0;	green_platform_transparency_texture[23][52] = 0;	green_platform_transparency_texture[23][53] = 0;	green_platform_transparency_texture[23][54] = 0;	green_platform_transparency_texture[23][55] = 0;	green_platform_transparency_texture[23][56] = 0;	green_platform_transparency_texture[23][57] = 0;	green_platform_transparency_texture[23][58] = 0;	green_platform_transparency_texture[23][59] = 0;	green_platform_transparency_texture[23][60] = 0;	green_platform_transparency_texture[23][61] = 0;	green_platform_transparency_texture[23][62] = 0;	green_platform_transparency_texture[23][63] = 0;	green_platform_transparency_texture[23][64] = 0;	green_platform_transparency_texture[23][65] = 0;	green_platform_transparency_texture[23][66] = 0;	green_platform_transparency_texture[23][67] = 0;	green_platform_transparency_texture[23][68] = 0;	green_platform_transparency_texture[23][69] = 0;	green_platform_transparency_texture[23][70] = 0;	green_platform_transparency_texture[23][71] = 0;	green_platform_transparency_texture[23][72] = 0;	green_platform_transparency_texture[23][73] = 0;	green_platform_transparency_texture[23][74] = 0;	green_platform_transparency_texture[23][75] = 0;	green_platform_transparency_texture[23][76] = 0;	green_platform_transparency_texture[23][77] = 0;	green_platform_transparency_texture[23][78] = 0;	green_platform_transparency_texture[23][79] = 0;	green_platform_transparency_texture[23][80] = 0;	green_platform_transparency_texture[23][81] = 0;	green_platform_transparency_texture[23][82] = 0;	green_platform_transparency_texture[23][83] = 0;	green_platform_transparency_texture[23][84] = 0;	green_platform_transparency_texture[23][85] = 0;	green_platform_transparency_texture[23][86] = 0;	green_platform_transparency_texture[23][87] = 0;	green_platform_transparency_texture[23][88] = 0;	green_platform_transparency_texture[23][89] = 0;	green_platform_transparency_texture[23][90] = 1;	green_platform_transparency_texture[23][91] = 1;	green_platform_transparency_texture[23][92] = 1;	green_platform_transparency_texture[23][93] = 1;	green_platform_transparency_texture[23][94] = 1;	green_platform_transparency_texture[23][95] = 1;	green_platform_transparency_texture[23][96] = 1;	green_platform_transparency_texture[23][97] = 1;	green_platform_transparency_texture[23][98] = 1;	green_platform_transparency_texture[23][99] = 1;	green_platform_transparency_texture[24][0] = 1;	green_platform_transparency_texture[24][1] = 1;	green_platform_transparency_texture[24][2] = 1;	green_platform_transparency_texture[24][3] = 1;	green_platform_transparency_texture[24][4] = 1;	green_platform_transparency_texture[24][5] = 1;	green_platform_transparency_texture[24][6] = 1;	green_platform_transparency_texture[24][7] = 1;	green_platform_transparency_texture[24][8] = 1;	green_platform_transparency_texture[24][9] = 0;	green_platform_transparency_texture[24][10] = 0;	green_platform_transparency_texture[24][11] = 0;	green_platform_transparency_texture[24][12] = 0;	green_platform_transparency_texture[24][13] = 0;	green_platform_transparency_texture[24][14] = 0;	green_platform_transparency_texture[24][15] = 0;	green_platform_transparency_texture[24][16] = 0;	green_platform_transparency_texture[24][17] = 0;	green_platform_transparency_texture[24][18] = 0;	green_platform_transparency_texture[24][19] = 0;	green_platform_transparency_texture[24][20] = 0;	green_platform_transparency_texture[24][21] = 0;	green_platform_transparency_texture[24][22] = 0;	green_platform_transparency_texture[24][23] = 0;	green_platform_transparency_texture[24][24] = 0;	green_platform_transparency_texture[24][25] = 0;	green_platform_transparency_texture[24][26] = 0;	green_platform_transparency_texture[24][27] = 0;	green_platform_transparency_texture[24][28] = 0;	green_platform_transparency_texture[24][29] = 0;	green_platform_transparency_texture[24][30] = 0;	green_platform_transparency_texture[24][31] = 0;	green_platform_transparency_texture[24][32] = 0;	green_platform_transparency_texture[24][33] = 0;	green_platform_transparency_texture[24][34] = 0;	green_platform_transparency_texture[24][35] = 0;	green_platform_transparency_texture[24][36] = 0;	green_platform_transparency_texture[24][37] = 0;	green_platform_transparency_texture[24][38] = 0;	green_platform_transparency_texture[24][39] = 0;	green_platform_transparency_texture[24][40] = 0;	green_platform_transparency_texture[24][41] = 0;	green_platform_transparency_texture[24][42] = 0;	green_platform_transparency_texture[24][43] = 0;	green_platform_transparency_texture[24][44] = 0;	green_platform_transparency_texture[24][45] = 0;	green_platform_transparency_texture[24][46] = 0;	green_platform_transparency_texture[24][47] = 0;	green_platform_transparency_texture[24][48] = 0;	green_platform_transparency_texture[24][49] = 0;	green_platform_transparency_texture[24][50] = 0;	green_platform_transparency_texture[24][51] = 0;	green_platform_transparency_texture[24][52] = 0;	green_platform_transparency_texture[24][53] = 0;	green_platform_transparency_texture[24][54] = 0;	green_platform_transparency_texture[24][55] = 0;	green_platform_transparency_texture[24][56] = 0;	green_platform_transparency_texture[24][57] = 0;	green_platform_transparency_texture[24][58] = 0;	green_platform_transparency_texture[24][59] = 0;	green_platform_transparency_texture[24][60] = 0;	green_platform_transparency_texture[24][61] = 0;	green_platform_transparency_texture[24][62] = 0;	green_platform_transparency_texture[24][63] = 0;	green_platform_transparency_texture[24][64] = 0;	green_platform_transparency_texture[24][65] = 0;	green_platform_transparency_texture[24][66] = 0;	green_platform_transparency_texture[24][67] = 0;	green_platform_transparency_texture[24][68] = 0;	green_platform_transparency_texture[24][69] = 0;	green_platform_transparency_texture[24][70] = 0;	green_platform_transparency_texture[24][71] = 0;	green_platform_transparency_texture[24][72] = 0;	green_platform_transparency_texture[24][73] = 0;	green_platform_transparency_texture[24][74] = 0;	green_platform_transparency_texture[24][75] = 0;	green_platform_transparency_texture[24][76] = 0;	green_platform_transparency_texture[24][77] = 0;	green_platform_transparency_texture[24][78] = 0;	green_platform_transparency_texture[24][79] = 0;	green_platform_transparency_texture[24][80] = 0;	green_platform_transparency_texture[24][81] = 0;	green_platform_transparency_texture[24][82] = 0;	green_platform_transparency_texture[24][83] = 0;	green_platform_transparency_texture[24][84] = 0;	green_platform_transparency_texture[24][85] = 0;	green_platform_transparency_texture[24][86] = 0;	green_platform_transparency_texture[24][87] = 0;	green_platform_transparency_texture[24][88] = 0;	green_platform_transparency_texture[24][89] = 0;	green_platform_transparency_texture[24][90] = 1;	green_platform_transparency_texture[24][91] = 1;	green_platform_transparency_texture[24][92] = 1;	green_platform_transparency_texture[24][93] = 1;	green_platform_transparency_texture[24][94] = 1;	green_platform_transparency_texture[24][95] = 1;	green_platform_transparency_texture[24][96] = 1;	green_platform_transparency_texture[24][97] = 1;	green_platform_transparency_texture[24][98] = 1;	green_platform_transparency_texture[24][99] = 1;	green_platform_transparency_texture[25][0] = 1;	green_platform_transparency_texture[25][1] = 1;	green_platform_transparency_texture[25][2] = 1;	green_platform_transparency_texture[25][3] = 1;	green_platform_transparency_texture[25][4] = 1;	green_platform_transparency_texture[25][5] = 1;	green_platform_transparency_texture[25][6] = 1;	green_platform_transparency_texture[25][7] = 1;	green_platform_transparency_texture[25][8] = 1;	green_platform_transparency_texture[25][9] = 1;	green_platform_transparency_texture[25][10] = 1;	green_platform_transparency_texture[25][11] = 1;	green_platform_transparency_texture[25][12] = 1;	green_platform_transparency_texture[25][13] = 1;	green_platform_transparency_texture[25][14] = 1;	green_platform_transparency_texture[25][15] = 1;	green_platform_transparency_texture[25][16] = 1;	green_platform_transparency_texture[25][17] = 1;	green_platform_transparency_texture[25][18] = 1;	green_platform_transparency_texture[25][19] = 1;	green_platform_transparency_texture[25][20] = 1;	green_platform_transparency_texture[25][21] = 1;	green_platform_transparency_texture[25][22] = 1;	green_platform_transparency_texture[25][23] = 1;	green_platform_transparency_texture[25][24] = 1;	green_platform_transparency_texture[25][25] = 1;	green_platform_transparency_texture[25][26] = 1;	green_platform_transparency_texture[25][27] = 1;	green_platform_transparency_texture[25][28] = 1;	green_platform_transparency_texture[25][29] = 1;	green_platform_transparency_texture[25][30] = 1;	green_platform_transparency_texture[25][31] = 1;	green_platform_transparency_texture[25][32] = 1;	green_platform_transparency_texture[25][33] = 1;	green_platform_transparency_texture[25][34] = 1;	green_platform_transparency_texture[25][35] = 1;	green_platform_transparency_texture[25][36] = 1;	green_platform_transparency_texture[25][37] = 1;	green_platform_transparency_texture[25][38] = 1;	green_platform_transparency_texture[25][39] = 1;	green_platform_transparency_texture[25][40] = 1;	green_platform_transparency_texture[25][41] = 1;	green_platform_transparency_texture[25][42] = 1;	green_platform_transparency_texture[25][43] = 1;	green_platform_transparency_texture[25][44] = 1;	green_platform_transparency_texture[25][45] = 1;	green_platform_transparency_texture[25][46] = 1;	green_platform_transparency_texture[25][47] = 1;	green_platform_transparency_texture[25][48] = 1;	green_platform_transparency_texture[25][49] = 1;	green_platform_transparency_texture[25][50] = 1;	green_platform_transparency_texture[25][51] = 1;	green_platform_transparency_texture[25][52] = 1;	green_platform_transparency_texture[25][53] = 1;	green_platform_transparency_texture[25][54] = 1;	green_platform_transparency_texture[25][55] = 1;	green_platform_transparency_texture[25][56] = 1;	green_platform_transparency_texture[25][57] = 1;	green_platform_transparency_texture[25][58] = 1;	green_platform_transparency_texture[25][59] = 1;	green_platform_transparency_texture[25][60] = 1;	green_platform_transparency_texture[25][61] = 1;	green_platform_transparency_texture[25][62] = 1;	green_platform_transparency_texture[25][63] = 1;	green_platform_transparency_texture[25][64] = 1;	green_platform_transparency_texture[25][65] = 1;	green_platform_transparency_texture[25][66] = 1;	green_platform_transparency_texture[25][67] = 1;	green_platform_transparency_texture[25][68] = 1;	green_platform_transparency_texture[25][69] = 1;	green_platform_transparency_texture[25][70] = 1;	green_platform_transparency_texture[25][71] = 1;	green_platform_transparency_texture[25][72] = 1;	green_platform_transparency_texture[25][73] = 1;	green_platform_transparency_texture[25][74] = 1;	green_platform_transparency_texture[25][75] = 1;	green_platform_transparency_texture[25][76] = 1;	green_platform_transparency_texture[25][77] = 1;	green_platform_transparency_texture[25][78] = 1;	green_platform_transparency_texture[25][79] = 1;	green_platform_transparency_texture[25][80] = 1;	green_platform_transparency_texture[25][81] = 1;	green_platform_transparency_texture[25][82] = 1;	green_platform_transparency_texture[25][83] = 1;	green_platform_transparency_texture[25][84] = 1;	green_platform_transparency_texture[25][85] = 1;	green_platform_transparency_texture[25][86] = 1;	green_platform_transparency_texture[25][87] = 1;	green_platform_transparency_texture[25][88] = 1;	green_platform_transparency_texture[25][89] = 1;	green_platform_transparency_texture[25][90] = 1;	green_platform_transparency_texture[25][91] = 1;	green_platform_transparency_texture[25][92] = 1;	green_platform_transparency_texture[25][93] = 1;	green_platform_transparency_texture[25][94] = 1;	green_platform_transparency_texture[25][95] = 1;	green_platform_transparency_texture[25][96] = 1;	green_platform_transparency_texture[25][97] = 1;	green_platform_transparency_texture[25][98] = 1;	green_platform_transparency_texture[25][99] = 1;	green_platform_transparency_texture[26][0] = 1;	green_platform_transparency_texture[26][1] = 1;	green_platform_transparency_texture[26][2] = 1;	green_platform_transparency_texture[26][3] = 1;	green_platform_transparency_texture[26][4] = 1;	green_platform_transparency_texture[26][5] = 1;	green_platform_transparency_texture[26][6] = 1;	green_platform_transparency_texture[26][7] = 1;	green_platform_transparency_texture[26][8] = 1;	green_platform_transparency_texture[26][9] = 1;	green_platform_transparency_texture[26][10] = 1;	green_platform_transparency_texture[26][11] = 1;	green_platform_transparency_texture[26][12] = 1;	green_platform_transparency_texture[26][13] = 1;	green_platform_transparency_texture[26][14] = 1;	green_platform_transparency_texture[26][15] = 1;	green_platform_transparency_texture[26][16] = 1;	green_platform_transparency_texture[26][17] = 1;	green_platform_transparency_texture[26][18] = 1;	green_platform_transparency_texture[26][19] = 1;	green_platform_transparency_texture[26][20] = 1;	green_platform_transparency_texture[26][21] = 1;	green_platform_transparency_texture[26][22] = 1;	green_platform_transparency_texture[26][23] = 1;	green_platform_transparency_texture[26][24] = 1;	green_platform_transparency_texture[26][25] = 1;	green_platform_transparency_texture[26][26] = 1;	green_platform_transparency_texture[26][27] = 1;	green_platform_transparency_texture[26][28] = 1;	green_platform_transparency_texture[26][29] = 1;	green_platform_transparency_texture[26][30] = 1;	green_platform_transparency_texture[26][31] = 1;	green_platform_transparency_texture[26][32] = 1;	green_platform_transparency_texture[26][33] = 1;	green_platform_transparency_texture[26][34] = 1;	green_platform_transparency_texture[26][35] = 1;	green_platform_transparency_texture[26][36] = 1;	green_platform_transparency_texture[26][37] = 1;	green_platform_transparency_texture[26][38] = 1;	green_platform_transparency_texture[26][39] = 1;	green_platform_transparency_texture[26][40] = 1;	green_platform_transparency_texture[26][41] = 1;	green_platform_transparency_texture[26][42] = 1;	green_platform_transparency_texture[26][43] = 1;	green_platform_transparency_texture[26][44] = 1;	green_platform_transparency_texture[26][45] = 1;	green_platform_transparency_texture[26][46] = 1;	green_platform_transparency_texture[26][47] = 1;	green_platform_transparency_texture[26][48] = 1;	green_platform_transparency_texture[26][49] = 1;	green_platform_transparency_texture[26][50] = 1;	green_platform_transparency_texture[26][51] = 1;	green_platform_transparency_texture[26][52] = 1;	green_platform_transparency_texture[26][53] = 1;	green_platform_transparency_texture[26][54] = 1;	green_platform_transparency_texture[26][55] = 1;	green_platform_transparency_texture[26][56] = 1;	green_platform_transparency_texture[26][57] = 1;	green_platform_transparency_texture[26][58] = 1;	green_platform_transparency_texture[26][59] = 1;	green_platform_transparency_texture[26][60] = 1;	green_platform_transparency_texture[26][61] = 1;	green_platform_transparency_texture[26][62] = 1;	green_platform_transparency_texture[26][63] = 1;	green_platform_transparency_texture[26][64] = 1;	green_platform_transparency_texture[26][65] = 1;	green_platform_transparency_texture[26][66] = 1;	green_platform_transparency_texture[26][67] = 1;	green_platform_transparency_texture[26][68] = 1;	green_platform_transparency_texture[26][69] = 1;	green_platform_transparency_texture[26][70] = 1;	green_platform_transparency_texture[26][71] = 1;	green_platform_transparency_texture[26][72] = 1;	green_platform_transparency_texture[26][73] = 1;	green_platform_transparency_texture[26][74] = 1;	green_platform_transparency_texture[26][75] = 1;	green_platform_transparency_texture[26][76] = 1;	green_platform_transparency_texture[26][77] = 1;	green_platform_transparency_texture[26][78] = 1;	green_platform_transparency_texture[26][79] = 1;	green_platform_transparency_texture[26][80] = 1;	green_platform_transparency_texture[26][81] = 1;	green_platform_transparency_texture[26][82] = 1;	green_platform_transparency_texture[26][83] = 1;	green_platform_transparency_texture[26][84] = 1;	green_platform_transparency_texture[26][85] = 1;	green_platform_transparency_texture[26][86] = 1;	green_platform_transparency_texture[26][87] = 1;	green_platform_transparency_texture[26][88] = 1;	green_platform_transparency_texture[26][89] = 1;	green_platform_transparency_texture[26][90] = 1;	green_platform_transparency_texture[26][91] = 1;	green_platform_transparency_texture[26][92] = 1;	green_platform_transparency_texture[26][93] = 1;	green_platform_transparency_texture[26][94] = 1;	green_platform_transparency_texture[26][95] = 1;	green_platform_transparency_texture[26][96] = 1;	green_platform_transparency_texture[26][97] = 1;	green_platform_transparency_texture[26][98] = 1;	green_platform_transparency_texture[26][99] = 1;	green_platform_transparency_texture[27][0] = 1;	green_platform_transparency_texture[27][1] = 1;	green_platform_transparency_texture[27][2] = 1;	green_platform_transparency_texture[27][3] = 1;	green_platform_transparency_texture[27][4] = 1;	green_platform_transparency_texture[27][5] = 1;	green_platform_transparency_texture[27][6] = 1;	green_platform_transparency_texture[27][7] = 1;	green_platform_transparency_texture[27][8] = 1;	green_platform_transparency_texture[27][9] = 1;	green_platform_transparency_texture[27][10] = 1;	green_platform_transparency_texture[27][11] = 1;	green_platform_transparency_texture[27][12] = 1;	green_platform_transparency_texture[27][13] = 1;	green_platform_transparency_texture[27][14] = 1;	green_platform_transparency_texture[27][15] = 1;	green_platform_transparency_texture[27][16] = 1;	green_platform_transparency_texture[27][17] = 1;	green_platform_transparency_texture[27][18] = 1;	green_platform_transparency_texture[27][19] = 1;	green_platform_transparency_texture[27][20] = 1;	green_platform_transparency_texture[27][21] = 1;	green_platform_transparency_texture[27][22] = 1;	green_platform_transparency_texture[27][23] = 1;	green_platform_transparency_texture[27][24] = 1;	green_platform_transparency_texture[27][25] = 1;	green_platform_transparency_texture[27][26] = 1;	green_platform_transparency_texture[27][27] = 1;	green_platform_transparency_texture[27][28] = 1;	green_platform_transparency_texture[27][29] = 1;	green_platform_transparency_texture[27][30] = 1;	green_platform_transparency_texture[27][31] = 1;	green_platform_transparency_texture[27][32] = 1;	green_platform_transparency_texture[27][33] = 1;	green_platform_transparency_texture[27][34] = 1;	green_platform_transparency_texture[27][35] = 1;	green_platform_transparency_texture[27][36] = 1;	green_platform_transparency_texture[27][37] = 1;	green_platform_transparency_texture[27][38] = 1;	green_platform_transparency_texture[27][39] = 1;	green_platform_transparency_texture[27][40] = 1;	green_platform_transparency_texture[27][41] = 1;	green_platform_transparency_texture[27][42] = 1;	green_platform_transparency_texture[27][43] = 1;	green_platform_transparency_texture[27][44] = 1;	green_platform_transparency_texture[27][45] = 1;	green_platform_transparency_texture[27][46] = 1;	green_platform_transparency_texture[27][47] = 1;	green_platform_transparency_texture[27][48] = 1;	green_platform_transparency_texture[27][49] = 1;	green_platform_transparency_texture[27][50] = 1;	green_platform_transparency_texture[27][51] = 1;	green_platform_transparency_texture[27][52] = 1;	green_platform_transparency_texture[27][53] = 1;	green_platform_transparency_texture[27][54] = 1;	green_platform_transparency_texture[27][55] = 1;	green_platform_transparency_texture[27][56] = 1;	green_platform_transparency_texture[27][57] = 1;	green_platform_transparency_texture[27][58] = 1;	green_platform_transparency_texture[27][59] = 1;	green_platform_transparency_texture[27][60] = 1;	green_platform_transparency_texture[27][61] = 1;	green_platform_transparency_texture[27][62] = 1;	green_platform_transparency_texture[27][63] = 1;	green_platform_transparency_texture[27][64] = 1;	green_platform_transparency_texture[27][65] = 1;	green_platform_transparency_texture[27][66] = 1;	green_platform_transparency_texture[27][67] = 1;	green_platform_transparency_texture[27][68] = 1;	green_platform_transparency_texture[27][69] = 1;	green_platform_transparency_texture[27][70] = 1;	green_platform_transparency_texture[27][71] = 1;	green_platform_transparency_texture[27][72] = 1;	green_platform_transparency_texture[27][73] = 1;	green_platform_transparency_texture[27][74] = 1;	green_platform_transparency_texture[27][75] = 1;	green_platform_transparency_texture[27][76] = 1;	green_platform_transparency_texture[27][77] = 1;	green_platform_transparency_texture[27][78] = 1;	green_platform_transparency_texture[27][79] = 1;	green_platform_transparency_texture[27][80] = 1;	green_platform_transparency_texture[27][81] = 1;	green_platform_transparency_texture[27][82] = 1;	green_platform_transparency_texture[27][83] = 1;	green_platform_transparency_texture[27][84] = 1;	green_platform_transparency_texture[27][85] = 1;	green_platform_transparency_texture[27][86] = 1;	green_platform_transparency_texture[27][87] = 1;	green_platform_transparency_texture[27][88] = 1;	green_platform_transparency_texture[27][89] = 1;	green_platform_transparency_texture[27][90] = 1;	green_platform_transparency_texture[27][91] = 1;	green_platform_transparency_texture[27][92] = 1;	green_platform_transparency_texture[27][93] = 1;	green_platform_transparency_texture[27][94] = 1;	green_platform_transparency_texture[27][95] = 1;	green_platform_transparency_texture[27][96] = 1;	green_platform_transparency_texture[27][97] = 1;	green_platform_transparency_texture[27][98] = 1;	green_platform_transparency_texture[27][99] = 1;	green_platform_transparency_texture[28][0] = 1;	green_platform_transparency_texture[28][1] = 1;	green_platform_transparency_texture[28][2] = 1;	green_platform_transparency_texture[28][3] = 1;	green_platform_transparency_texture[28][4] = 1;	green_platform_transparency_texture[28][5] = 1;	green_platform_transparency_texture[28][6] = 1;	green_platform_transparency_texture[28][7] = 1;	green_platform_transparency_texture[28][8] = 1;	green_platform_transparency_texture[28][9] = 1;	green_platform_transparency_texture[28][10] = 1;	green_platform_transparency_texture[28][11] = 1;	green_platform_transparency_texture[28][12] = 1;	green_platform_transparency_texture[28][13] = 1;	green_platform_transparency_texture[28][14] = 1;	green_platform_transparency_texture[28][15] = 1;	green_platform_transparency_texture[28][16] = 1;	green_platform_transparency_texture[28][17] = 1;	green_platform_transparency_texture[28][18] = 1;	green_platform_transparency_texture[28][19] = 1;	green_platform_transparency_texture[28][20] = 1;	green_platform_transparency_texture[28][21] = 1;	green_platform_transparency_texture[28][22] = 1;	green_platform_transparency_texture[28][23] = 1;	green_platform_transparency_texture[28][24] = 1;	green_platform_transparency_texture[28][25] = 1;	green_platform_transparency_texture[28][26] = 1;	green_platform_transparency_texture[28][27] = 1;	green_platform_transparency_texture[28][28] = 1;	green_platform_transparency_texture[28][29] = 1;	green_platform_transparency_texture[28][30] = 1;	green_platform_transparency_texture[28][31] = 1;	green_platform_transparency_texture[28][32] = 1;	green_platform_transparency_texture[28][33] = 1;	green_platform_transparency_texture[28][34] = 1;	green_platform_transparency_texture[28][35] = 1;	green_platform_transparency_texture[28][36] = 1;	green_platform_transparency_texture[28][37] = 1;	green_platform_transparency_texture[28][38] = 1;	green_platform_transparency_texture[28][39] = 1;	green_platform_transparency_texture[28][40] = 1;	green_platform_transparency_texture[28][41] = 1;	green_platform_transparency_texture[28][42] = 1;	green_platform_transparency_texture[28][43] = 1;	green_platform_transparency_texture[28][44] = 1;	green_platform_transparency_texture[28][45] = 1;	green_platform_transparency_texture[28][46] = 1;	green_platform_transparency_texture[28][47] = 1;	green_platform_transparency_texture[28][48] = 1;	green_platform_transparency_texture[28][49] = 1;	green_platform_transparency_texture[28][50] = 1;	green_platform_transparency_texture[28][51] = 1;	green_platform_transparency_texture[28][52] = 1;	green_platform_transparency_texture[28][53] = 1;	green_platform_transparency_texture[28][54] = 1;	green_platform_transparency_texture[28][55] = 1;	green_platform_transparency_texture[28][56] = 1;	green_platform_transparency_texture[28][57] = 1;	green_platform_transparency_texture[28][58] = 1;	green_platform_transparency_texture[28][59] = 1;	green_platform_transparency_texture[28][60] = 1;	green_platform_transparency_texture[28][61] = 1;	green_platform_transparency_texture[28][62] = 1;	green_platform_transparency_texture[28][63] = 1;	green_platform_transparency_texture[28][64] = 1;	green_platform_transparency_texture[28][65] = 1;	green_platform_transparency_texture[28][66] = 1;	green_platform_transparency_texture[28][67] = 1;	green_platform_transparency_texture[28][68] = 1;	green_platform_transparency_texture[28][69] = 1;	green_platform_transparency_texture[28][70] = 1;	green_platform_transparency_texture[28][71] = 1;	green_platform_transparency_texture[28][72] = 1;	green_platform_transparency_texture[28][73] = 1;	green_platform_transparency_texture[28][74] = 1;	green_platform_transparency_texture[28][75] = 1;	green_platform_transparency_texture[28][76] = 1;	green_platform_transparency_texture[28][77] = 1;	green_platform_transparency_texture[28][78] = 1;	green_platform_transparency_texture[28][79] = 1;	green_platform_transparency_texture[28][80] = 1;	green_platform_transparency_texture[28][81] = 1;	green_platform_transparency_texture[28][82] = 1;	green_platform_transparency_texture[28][83] = 1;	green_platform_transparency_texture[28][84] = 1;	green_platform_transparency_texture[28][85] = 1;	green_platform_transparency_texture[28][86] = 1;	green_platform_transparency_texture[28][87] = 1;	green_platform_transparency_texture[28][88] = 1;	green_platform_transparency_texture[28][89] = 1;	green_platform_transparency_texture[28][90] = 1;	green_platform_transparency_texture[28][91] = 1;	green_platform_transparency_texture[28][92] = 1;	green_platform_transparency_texture[28][93] = 1;	green_platform_transparency_texture[28][94] = 1;	green_platform_transparency_texture[28][95] = 1;	green_platform_transparency_texture[28][96] = 1;	green_platform_transparency_texture[28][97] = 1;	green_platform_transparency_texture[28][98] = 1;	green_platform_transparency_texture[28][99] = 1;	green_platform_transparency_texture[29][0] = 1;	green_platform_transparency_texture[29][1] = 1;	green_platform_transparency_texture[29][2] = 1;	green_platform_transparency_texture[29][3] = 1;	green_platform_transparency_texture[29][4] = 1;	green_platform_transparency_texture[29][5] = 1;	green_platform_transparency_texture[29][6] = 1;	green_platform_transparency_texture[29][7] = 1;	green_platform_transparency_texture[29][8] = 1;	green_platform_transparency_texture[29][9] = 1;	green_platform_transparency_texture[29][10] = 1;	green_platform_transparency_texture[29][11] = 1;	green_platform_transparency_texture[29][12] = 1;	green_platform_transparency_texture[29][13] = 1;	green_platform_transparency_texture[29][14] = 1;	green_platform_transparency_texture[29][15] = 1;	green_platform_transparency_texture[29][16] = 1;	green_platform_transparency_texture[29][17] = 1;	green_platform_transparency_texture[29][18] = 1;	green_platform_transparency_texture[29][19] = 1;	green_platform_transparency_texture[29][20] = 1;	green_platform_transparency_texture[29][21] = 1;	green_platform_transparency_texture[29][22] = 1;	green_platform_transparency_texture[29][23] = 1;	green_platform_transparency_texture[29][24] = 1;	green_platform_transparency_texture[29][25] = 1;	green_platform_transparency_texture[29][26] = 1;	green_platform_transparency_texture[29][27] = 1;	green_platform_transparency_texture[29][28] = 1;	green_platform_transparency_texture[29][29] = 1;	green_platform_transparency_texture[29][30] = 1;	green_platform_transparency_texture[29][31] = 1;	green_platform_transparency_texture[29][32] = 1;	green_platform_transparency_texture[29][33] = 1;	green_platform_transparency_texture[29][34] = 1;	green_platform_transparency_texture[29][35] = 1;	green_platform_transparency_texture[29][36] = 1;	green_platform_transparency_texture[29][37] = 1;	green_platform_transparency_texture[29][38] = 1;	green_platform_transparency_texture[29][39] = 1;	green_platform_transparency_texture[29][40] = 1;	green_platform_transparency_texture[29][41] = 1;	green_platform_transparency_texture[29][42] = 1;	green_platform_transparency_texture[29][43] = 1;	green_platform_transparency_texture[29][44] = 1;	green_platform_transparency_texture[29][45] = 1;	green_platform_transparency_texture[29][46] = 1;	green_platform_transparency_texture[29][47] = 1;	green_platform_transparency_texture[29][48] = 1;	green_platform_transparency_texture[29][49] = 1;	green_platform_transparency_texture[29][50] = 1;	green_platform_transparency_texture[29][51] = 1;	green_platform_transparency_texture[29][52] = 1;	green_platform_transparency_texture[29][53] = 1;	green_platform_transparency_texture[29][54] = 1;	green_platform_transparency_texture[29][55] = 1;	green_platform_transparency_texture[29][56] = 1;	green_platform_transparency_texture[29][57] = 1;	green_platform_transparency_texture[29][58] = 1;	green_platform_transparency_texture[29][59] = 1;	green_platform_transparency_texture[29][60] = 1;	green_platform_transparency_texture[29][61] = 1;	green_platform_transparency_texture[29][62] = 1;	green_platform_transparency_texture[29][63] = 1;	green_platform_transparency_texture[29][64] = 1;	green_platform_transparency_texture[29][65] = 1;	green_platform_transparency_texture[29][66] = 1;	green_platform_transparency_texture[29][67] = 1;	green_platform_transparency_texture[29][68] = 1;	green_platform_transparency_texture[29][69] = 1;	green_platform_transparency_texture[29][70] = 1;	green_platform_transparency_texture[29][71] = 1;	green_platform_transparency_texture[29][72] = 1;	green_platform_transparency_texture[29][73] = 1;	green_platform_transparency_texture[29][74] = 1;	green_platform_transparency_texture[29][75] = 1;	green_platform_transparency_texture[29][76] = 1;	green_platform_transparency_texture[29][77] = 1;	green_platform_transparency_texture[29][78] = 1;	green_platform_transparency_texture[29][79] = 1;	green_platform_transparency_texture[29][80] = 1;	green_platform_transparency_texture[29][81] = 1;	green_platform_transparency_texture[29][82] = 1;	green_platform_transparency_texture[29][83] = 1;	green_platform_transparency_texture[29][84] = 1;	green_platform_transparency_texture[29][85] = 1;	green_platform_transparency_texture[29][86] = 1;	green_platform_transparency_texture[29][87] = 1;	green_platform_transparency_texture[29][88] = 1;	green_platform_transparency_texture[29][89] = 1;	green_platform_transparency_texture[29][90] = 1;	green_platform_transparency_texture[29][91] = 1;	green_platform_transparency_texture[29][92] = 1;	green_platform_transparency_texture[29][93] = 1;	green_platform_transparency_texture[29][94] = 1;	green_platform_transparency_texture[29][95] = 1;	green_platform_transparency_texture[29][96] = 1;	green_platform_transparency_texture[29][97] = 1;	green_platform_transparency_texture[29][98] = 1;	green_platform_transparency_texture[29][99] = 1;
end

endmodule
