module platforms(
	output [4:0][3:0][:] platforms
)



endmodule
