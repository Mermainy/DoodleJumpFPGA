`ifndef INITIAL_FOUR_TRANSPARENT

// Module definition:
// logic [11:0][12:0][2:0][3:0] four_transparent_rgb;
// logic [11:0][12:0] four_transparent_alpha;

`define INITIAL_FOUR_TRANSPARENT \
always_comb begin \
	four_transparent_rgb[0][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][2] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][3] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][4] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][5] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][6] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][7] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[0][8] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[0][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[0][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[0][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[0][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][2] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][3] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][4] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][5] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][6] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[1][7] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[1][8] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[1][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[1][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[1][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[1][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[2][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[2][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[2][2] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[2][3] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[2][4] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[2][5] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[2][6] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[2][7] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[2][8] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[2][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[2][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[2][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[2][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[3][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[3][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[3][2] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[3][3] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[3][4] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[3][5] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[3][6] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[3][7] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[3][8] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[3][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[3][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[3][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[3][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[4][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[4][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[4][2] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[4][3] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[4][4] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[4][5] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[4][6] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[4][7] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[4][8] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[4][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[4][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[4][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[4][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[5][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[5][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[5][2] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[5][3] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[5][4] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[5][5] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[5][6] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[5][7] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[5][8] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[5][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[5][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[5][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[5][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[6][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[6][1] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[6][2] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[6][3] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[6][4] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[6][5] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[6][6] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[6][7] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[6][8] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[6][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[6][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[6][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[6][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[7][0] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[7][1] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[7][2] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[7][3] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[7][4] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[7][5] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[7][6] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[7][7] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[7][8] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[7][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[7][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[7][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[7][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[8][0] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][1] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][2] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][3] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][4] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][5] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][6] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][7] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][8] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[8][12] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][0] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][1] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][2] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][3] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][4] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][5] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][6] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][7] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][8] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[9][12] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[10][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][2] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][3] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][4] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][5] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][6] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][7] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][8] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[10][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[10][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[10][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[10][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][0] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][1] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][2] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][3] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][4] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][5] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][6] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][7] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][8] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_rgb[11][9] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[11][10] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[11][11] = {4'b0, 4'b0, 4'b0}; \
	four_transparent_rgb[11][12] = {4'b1111, 4'b1111, 4'b1111}; \
	four_transparent_alpha[0][0] = 1'b1; \
	four_transparent_alpha[0][1] = 1'b1; \
	four_transparent_alpha[0][2] = 1'b1; \
	four_transparent_alpha[0][3] = 1'b1; \
	four_transparent_alpha[0][4] = 1'b1; \
	four_transparent_alpha[0][5] = 1'b1; \
	four_transparent_alpha[0][6] = 1'b1; \
	four_transparent_alpha[0][7] = 1'b1; \
	four_transparent_alpha[0][8] = 1'b0; \
	four_transparent_alpha[0][9] = 1'b0; \
	four_transparent_alpha[0][10] = 1'b0; \
	four_transparent_alpha[0][11] = 1'b0; \
	four_transparent_alpha[0][12] = 1'b1; \
	four_transparent_alpha[1][0] = 1'b1; \
	four_transparent_alpha[1][1] = 1'b1; \
	four_transparent_alpha[1][2] = 1'b1; \
	four_transparent_alpha[1][3] = 1'b1; \
	four_transparent_alpha[1][4] = 1'b1; \
	four_transparent_alpha[1][5] = 1'b1; \
	four_transparent_alpha[1][6] = 1'b1; \
	four_transparent_alpha[1][7] = 1'b0; \
	four_transparent_alpha[1][8] = 1'b0; \
	four_transparent_alpha[1][9] = 1'b0; \
	four_transparent_alpha[1][10] = 1'b0; \
	four_transparent_alpha[1][11] = 1'b0; \
	four_transparent_alpha[1][12] = 1'b1; \
	four_transparent_alpha[2][0] = 1'b1; \
	four_transparent_alpha[2][1] = 1'b1; \
	four_transparent_alpha[2][2] = 1'b1; \
	four_transparent_alpha[2][3] = 1'b1; \
	four_transparent_alpha[2][4] = 1'b1; \
	four_transparent_alpha[2][5] = 1'b1; \
	four_transparent_alpha[2][6] = 1'b0; \
	four_transparent_alpha[2][7] = 1'b0; \
	four_transparent_alpha[2][8] = 1'b0; \
	four_transparent_alpha[2][9] = 1'b0; \
	four_transparent_alpha[2][10] = 1'b0; \
	four_transparent_alpha[2][11] = 1'b0; \
	four_transparent_alpha[2][12] = 1'b1; \
	four_transparent_alpha[3][0] = 1'b1; \
	four_transparent_alpha[3][1] = 1'b1; \
	four_transparent_alpha[3][2] = 1'b1; \
	four_transparent_alpha[3][3] = 1'b1; \
	four_transparent_alpha[3][4] = 1'b0; \
	four_transparent_alpha[3][5] = 1'b0; \
	four_transparent_alpha[3][6] = 1'b0; \
	four_transparent_alpha[3][7] = 1'b0; \
	four_transparent_alpha[3][8] = 1'b1; \
	four_transparent_alpha[3][9] = 1'b0; \
	four_transparent_alpha[3][10] = 1'b0; \
	four_transparent_alpha[3][11] = 1'b0; \
	four_transparent_alpha[3][12] = 1'b1; \
	four_transparent_alpha[4][0] = 1'b1; \
	four_transparent_alpha[4][1] = 1'b1; \
	four_transparent_alpha[4][2] = 1'b1; \
	four_transparent_alpha[4][3] = 1'b0; \
	four_transparent_alpha[4][4] = 1'b0; \
	four_transparent_alpha[4][5] = 1'b0; \
	four_transparent_alpha[4][6] = 1'b0; \
	four_transparent_alpha[4][7] = 1'b1; \
	four_transparent_alpha[4][8] = 1'b1; \
	four_transparent_alpha[4][9] = 1'b0; \
	four_transparent_alpha[4][10] = 1'b0; \
	four_transparent_alpha[4][11] = 1'b0; \
	four_transparent_alpha[4][12] = 1'b1; \
	four_transparent_alpha[5][0] = 1'b1; \
	four_transparent_alpha[5][1] = 1'b1; \
	four_transparent_alpha[5][2] = 1'b0; \
	four_transparent_alpha[5][3] = 1'b0; \
	four_transparent_alpha[5][4] = 1'b0; \
	four_transparent_alpha[5][5] = 1'b0; \
	four_transparent_alpha[5][6] = 1'b1; \
	four_transparent_alpha[5][7] = 1'b1; \
	four_transparent_alpha[5][8] = 1'b1; \
	four_transparent_alpha[5][9] = 1'b0; \
	four_transparent_alpha[5][10] = 1'b0; \
	four_transparent_alpha[5][11] = 1'b0; \
	four_transparent_alpha[5][12] = 1'b1; \
	four_transparent_alpha[6][0] = 1'b1; \
	four_transparent_alpha[6][1] = 1'b0; \
	four_transparent_alpha[6][2] = 1'b0; \
	four_transparent_alpha[6][3] = 1'b0; \
	four_transparent_alpha[6][4] = 1'b0; \
	four_transparent_alpha[6][5] = 1'b1; \
	four_transparent_alpha[6][6] = 1'b1; \
	four_transparent_alpha[6][7] = 1'b1; \
	four_transparent_alpha[6][8] = 1'b1; \
	four_transparent_alpha[6][9] = 1'b0; \
	four_transparent_alpha[6][10] = 1'b0; \
	four_transparent_alpha[6][11] = 1'b0; \
	four_transparent_alpha[6][12] = 1'b1; \
	four_transparent_alpha[7][0] = 1'b0; \
	four_transparent_alpha[7][1] = 1'b0; \
	four_transparent_alpha[7][2] = 1'b0; \
	four_transparent_alpha[7][3] = 1'b1; \
	four_transparent_alpha[7][4] = 1'b1; \
	four_transparent_alpha[7][5] = 1'b1; \
	four_transparent_alpha[7][6] = 1'b1; \
	four_transparent_alpha[7][7] = 1'b1; \
	four_transparent_alpha[7][8] = 1'b1; \
	four_transparent_alpha[7][9] = 1'b0; \
	four_transparent_alpha[7][10] = 1'b0; \
	four_transparent_alpha[7][11] = 1'b0; \
	four_transparent_alpha[7][12] = 1'b1; \
	four_transparent_alpha[8][0] = 1'b0; \
	four_transparent_alpha[8][1] = 1'b0; \
	four_transparent_alpha[8][2] = 1'b0; \
	four_transparent_alpha[8][3] = 1'b0; \
	four_transparent_alpha[8][4] = 1'b0; \
	four_transparent_alpha[8][5] = 1'b0; \
	four_transparent_alpha[8][6] = 1'b0; \
	four_transparent_alpha[8][7] = 1'b0; \
	four_transparent_alpha[8][8] = 1'b0; \
	four_transparent_alpha[8][9] = 1'b0; \
	four_transparent_alpha[8][10] = 1'b0; \
	four_transparent_alpha[8][11] = 1'b0; \
	four_transparent_alpha[8][12] = 1'b0; \
	four_transparent_alpha[9][0] = 1'b0; \
	four_transparent_alpha[9][1] = 1'b0; \
	four_transparent_alpha[9][2] = 1'b0; \
	four_transparent_alpha[9][3] = 1'b0; \
	four_transparent_alpha[9][4] = 1'b0; \
	four_transparent_alpha[9][5] = 1'b0; \
	four_transparent_alpha[9][6] = 1'b0; \
	four_transparent_alpha[9][7] = 1'b0; \
	four_transparent_alpha[9][8] = 1'b0; \
	four_transparent_alpha[9][9] = 1'b0; \
	four_transparent_alpha[9][10] = 1'b0; \
	four_transparent_alpha[9][11] = 1'b0; \
	four_transparent_alpha[9][12] = 1'b0; \
	four_transparent_alpha[10][0] = 1'b1; \
	four_transparent_alpha[10][1] = 1'b1; \
	four_transparent_alpha[10][2] = 1'b1; \
	four_transparent_alpha[10][3] = 1'b1; \
	four_transparent_alpha[10][4] = 1'b1; \
	four_transparent_alpha[10][5] = 1'b1; \
	four_transparent_alpha[10][6] = 1'b1; \
	four_transparent_alpha[10][7] = 1'b1; \
	four_transparent_alpha[10][8] = 1'b1; \
	four_transparent_alpha[10][9] = 1'b0; \
	four_transparent_alpha[10][10] = 1'b0; \
	four_transparent_alpha[10][11] = 1'b0; \
	four_transparent_alpha[10][12] = 1'b1; \
	four_transparent_alpha[11][0] = 1'b1; \
	four_transparent_alpha[11][1] = 1'b1; \
	four_transparent_alpha[11][2] = 1'b1; \
	four_transparent_alpha[11][3] = 1'b1; \
	four_transparent_alpha[11][4] = 1'b1; \
	four_transparent_alpha[11][5] = 1'b1; \
	four_transparent_alpha[11][6] = 1'b1; \
	four_transparent_alpha[11][7] = 1'b1; \
	four_transparent_alpha[11][8] = 1'b1; \
	four_transparent_alpha[11][9] = 1'b0; \
	four_transparent_alpha[11][10] = 1'b0; \
	four_transparent_alpha[11][11] = 1'b0; \
	four_transparent_alpha[11][12] = 1'b1; \
end

`endif // INITIAL_FOUR_TRANSPARENT
