module doodle # (
	parameter int unsigned VELOCITY = 44,
	parameter int unsigned ACCELERATION = 4,
	parameter int unsigned FPS = 50,
	parameter int unsigned CLK = 50000000
) (
	input clk,
	input rst,
	input [1:0][9:0] ground,
	
	input [10:0] beam_x,
	input [9:0] beam_y,
	
	input signed [8:0] delta_x,
	output logic [9:0] doodle_y,
	output logic signed [11:0] doodle_x,
	output logic [2:0][3:0] color,
	output logic is_transparent
);




logic [79:0][79:0][2:0][3:0] doodle_right_texture;
logic [79:0][79:0] doodle_right_transparency_texture;
logic [79:0][79:0][2:0][3:0] doodle_left_texture;
logic [79:0][79:0] doodle_left_transparency_texture;


logic draw;


assign draw = doodle_x <= beam_x && beam_x < doodle_x + 80 - 2 
		&& doodle_y <= beam_y && beam_y < doodle_y + 80 - 1;

logic previous_texture_direction;  // 1 - left
always_ff @ (posedge clk) begin
	if (rst) begin
		previous_texture_direction <= 0;
	end else begin
		if (draw) begin
			if (delta_x < 0 || delta_x == 0 && previous_texture_direction) begin
				previous_texture_direction = 1;
				color[0] = doodle_left_texture[beam_y - doodle_y][beam_x - doodle_x][0];
				color[1] = doodle_left_texture[beam_y - doodle_y][beam_x - doodle_x][1];
				color[2] = doodle_left_texture[beam_y - doodle_y][beam_x - doodle_x][2];
				is_transparent = doodle_left_transparency_texture[beam_y - doodle_y][beam_x - doodle_x];
			end else begin
				previous_texture_direction = 0;
				color[0] = doodle_right_texture[beam_y - doodle_y][beam_x - doodle_x][0];
				color[1] = doodle_right_texture[beam_y - doodle_y][beam_x - doodle_x][1];
				color[2] = doodle_right_texture[beam_y - doodle_y][beam_x - doodle_x][2];
				is_transparent = doodle_right_transparency_texture[beam_y - doodle_y][beam_x - doodle_x];
			end
		end else begin 
			is_transparent = 1; 
			previous_texture_direction = previous_texture_direction;
		end
	end
end

logic [$clog2(CLK / FPS):0] fps_counter; 
logic [7:0] jump_counter;
// position
always_ff @ (posedge clk) begin
	if (rst) begin
		doodle_x <= 472;
		doodle_y <= 688;
	end else begin
		fps_counter <= fps_counter + 1;
		if (&fps_counter) begin
			if (doodle_x <= 300) 
				doodle_x <= 641;
			else if (doodle_x >= 642) 
				doodle_x <= 301;
			else 
				doodle_x <= doodle_x + delta_x;
			
			if (doodle_y + 80 >= ground[0] && ground[1] <= doodle_x 
			&& doodle_x <= ground[0] + 100) begin
				doodle_y <= ground - 1;
				jump_counter <= 1;
			end else begin
				doodle_y <= ground - VELOCITY * jump_counter + ACCELERATION * jump_counter * jump_counter / 2;
				jump_counter <= jump_counter + 1;
			end
		end
	end
end


always_comb begin
		doodle_right_texture[0][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[0][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[1][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[2][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[3][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[4][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[5][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[6][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[7][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[8][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[9][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[10][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[11][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[12][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[12][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[13][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[13][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[14][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[14][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[15][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[15][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[16][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[16][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[17][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[17][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[18][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[18][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[19][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[19][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[20][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[20][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[21][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[21][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[22][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[22][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[23][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[23][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[24][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[24][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[25][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[25][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[26][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[26][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[27][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[27][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][52] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][53] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][54] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][55] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][56] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][57] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][58] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][59] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][60] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][61] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][62] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][63] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][68] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][69] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][70] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][71] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[28][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[28][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][52] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][53] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][54] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][55] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][56] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][57] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][58] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][59] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][60] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][61] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][62] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][63] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][68] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][69] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][70] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][71] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[29][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[29][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][52] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][53] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][54] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][55] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][56] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][57] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][58] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][59] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][60] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][61] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][62] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][63] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][68] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][69] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][70] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][71] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[30][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[30][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][52] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][53] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][54] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][55] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][56] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][57] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][58] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][59] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][60] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][61] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][62] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][63] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][68] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][69] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][70] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][71] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[31][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[31][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[32][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[32][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[33][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[33][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[34][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[34][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][48] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][49] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][50] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][51] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[35][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[35][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[36][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[36][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[37][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[37][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[38][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[38][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[39][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[39][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[40][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[40][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[41][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[41][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[42][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[42][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[43][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[43][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[44][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[45][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[46][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[47][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[48][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[48][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[49][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[49][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[50][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[50][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[51][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[51][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[52][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[52][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[53][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[53][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[54][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[54][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][8] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][9] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][10] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][11] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][12] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][13] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][14] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][15] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][16] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][17] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][18] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][19] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][20] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][21] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][22] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][23] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][24] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][25] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][26] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][27] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][28] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][29] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][30] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][31] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][32] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][33] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][34] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][35] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][36] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][37] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][38] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][39] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][40] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][41] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][42] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][43] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][44] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][45] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][46] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][47] = {4'b0, 4'b1111, 4'b0};	doodle_right_texture[55][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[55][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[56][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[57][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[58][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[59][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[60][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[61][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[62][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[63][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[64][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[65][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[66][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[67][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[68][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[69][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[70][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[71][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[72][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[73][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[74][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[75][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[76][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[77][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[78][79] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][0] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][1] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][2] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][3] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][4] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][5] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][6] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][7] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][8] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][9] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][10] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][11] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][12] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][13] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][14] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][15] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][16] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][17] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][18] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][19] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][20] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][21] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][22] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][23] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][24] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][25] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][26] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][27] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][28] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][29] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][30] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][31] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][32] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][33] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][34] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][35] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][36] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][37] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][38] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][39] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][40] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][41] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][42] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][43] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][44] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][45] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][46] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][47] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][48] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][49] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][50] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][51] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][52] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][53] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][54] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][55] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][56] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][57] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][58] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][59] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][60] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][61] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][62] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][63] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][64] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][65] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][66] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][67] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][68] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][69] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][70] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][71] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][72] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][73] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][74] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][75] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][76] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][77] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][78] = {4'b0, 4'b0, 4'b0};	doodle_right_texture[79][79] = {4'b0, 4'b0, 4'b0};
		doodle_right_transparency_texture[0][0] = 1;	doodle_right_transparency_texture[0][1] = 1;	doodle_right_transparency_texture[0][2] = 1;	doodle_right_transparency_texture[0][3] = 1;	doodle_right_transparency_texture[0][4] = 1;	doodle_right_transparency_texture[0][5] = 1;	doodle_right_transparency_texture[0][6] = 1;	doodle_right_transparency_texture[0][7] = 1;	doodle_right_transparency_texture[0][8] = 1;	doodle_right_transparency_texture[0][9] = 1;	doodle_right_transparency_texture[0][10] = 1;	doodle_right_transparency_texture[0][11] = 1;	doodle_right_transparency_texture[0][12] = 1;	doodle_right_transparency_texture[0][13] = 1;	doodle_right_transparency_texture[0][14] = 1;	doodle_right_transparency_texture[0][15] = 1;	doodle_right_transparency_texture[0][16] = 1;	doodle_right_transparency_texture[0][17] = 1;	doodle_right_transparency_texture[0][18] = 1;	doodle_right_transparency_texture[0][19] = 1;	doodle_right_transparency_texture[0][20] = 1;	doodle_right_transparency_texture[0][21] = 1;	doodle_right_transparency_texture[0][22] = 1;	doodle_right_transparency_texture[0][23] = 1;	doodle_right_transparency_texture[0][24] = 1;	doodle_right_transparency_texture[0][25] = 1;	doodle_right_transparency_texture[0][26] = 1;	doodle_right_transparency_texture[0][27] = 1;	doodle_right_transparency_texture[0][28] = 1;	doodle_right_transparency_texture[0][29] = 1;	doodle_right_transparency_texture[0][30] = 1;	doodle_right_transparency_texture[0][31] = 1;	doodle_right_transparency_texture[0][32] = 1;	doodle_right_transparency_texture[0][33] = 1;	doodle_right_transparency_texture[0][34] = 1;	doodle_right_transparency_texture[0][35] = 1;	doodle_right_transparency_texture[0][36] = 1;	doodle_right_transparency_texture[0][37] = 1;	doodle_right_transparency_texture[0][38] = 1;	doodle_right_transparency_texture[0][39] = 1;	doodle_right_transparency_texture[0][40] = 1;	doodle_right_transparency_texture[0][41] = 1;	doodle_right_transparency_texture[0][42] = 1;	doodle_right_transparency_texture[0][43] = 1;	doodle_right_transparency_texture[0][44] = 1;	doodle_right_transparency_texture[0][45] = 1;	doodle_right_transparency_texture[0][46] = 1;	doodle_right_transparency_texture[0][47] = 1;	doodle_right_transparency_texture[0][48] = 1;	doodle_right_transparency_texture[0][49] = 1;	doodle_right_transparency_texture[0][50] = 1;	doodle_right_transparency_texture[0][51] = 1;	doodle_right_transparency_texture[0][52] = 1;	doodle_right_transparency_texture[0][53] = 1;	doodle_right_transparency_texture[0][54] = 1;	doodle_right_transparency_texture[0][55] = 1;	doodle_right_transparency_texture[0][56] = 1;	doodle_right_transparency_texture[0][57] = 1;	doodle_right_transparency_texture[0][58] = 1;	doodle_right_transparency_texture[0][59] = 1;	doodle_right_transparency_texture[0][60] = 1;	doodle_right_transparency_texture[0][61] = 1;	doodle_right_transparency_texture[0][62] = 1;	doodle_right_transparency_texture[0][63] = 1;	doodle_right_transparency_texture[0][64] = 1;	doodle_right_transparency_texture[0][65] = 1;	doodle_right_transparency_texture[0][66] = 1;	doodle_right_transparency_texture[0][67] = 1;	doodle_right_transparency_texture[0][68] = 1;	doodle_right_transparency_texture[0][69] = 1;	doodle_right_transparency_texture[0][70] = 1;	doodle_right_transparency_texture[0][71] = 1;	doodle_right_transparency_texture[0][72] = 1;	doodle_right_transparency_texture[0][73] = 1;	doodle_right_transparency_texture[0][74] = 1;	doodle_right_transparency_texture[0][75] = 1;	doodle_right_transparency_texture[0][76] = 1;	doodle_right_transparency_texture[0][77] = 1;	doodle_right_transparency_texture[0][78] = 1;	doodle_right_transparency_texture[0][79] = 1;	doodle_right_transparency_texture[1][0] = 1;	doodle_right_transparency_texture[1][1] = 1;	doodle_right_transparency_texture[1][2] = 1;	doodle_right_transparency_texture[1][3] = 1;	doodle_right_transparency_texture[1][4] = 1;	doodle_right_transparency_texture[1][5] = 1;	doodle_right_transparency_texture[1][6] = 1;	doodle_right_transparency_texture[1][7] = 1;	doodle_right_transparency_texture[1][8] = 1;	doodle_right_transparency_texture[1][9] = 1;	doodle_right_transparency_texture[1][10] = 1;	doodle_right_transparency_texture[1][11] = 1;	doodle_right_transparency_texture[1][12] = 1;	doodle_right_transparency_texture[1][13] = 1;	doodle_right_transparency_texture[1][14] = 1;	doodle_right_transparency_texture[1][15] = 1;	doodle_right_transparency_texture[1][16] = 1;	doodle_right_transparency_texture[1][17] = 1;	doodle_right_transparency_texture[1][18] = 1;	doodle_right_transparency_texture[1][19] = 1;	doodle_right_transparency_texture[1][20] = 1;	doodle_right_transparency_texture[1][21] = 1;	doodle_right_transparency_texture[1][22] = 1;	doodle_right_transparency_texture[1][23] = 1;	doodle_right_transparency_texture[1][24] = 1;	doodle_right_transparency_texture[1][25] = 1;	doodle_right_transparency_texture[1][26] = 1;	doodle_right_transparency_texture[1][27] = 1;	doodle_right_transparency_texture[1][28] = 1;	doodle_right_transparency_texture[1][29] = 1;	doodle_right_transparency_texture[1][30] = 1;	doodle_right_transparency_texture[1][31] = 1;	doodle_right_transparency_texture[1][32] = 1;	doodle_right_transparency_texture[1][33] = 1;	doodle_right_transparency_texture[1][34] = 1;	doodle_right_transparency_texture[1][35] = 1;	doodle_right_transparency_texture[1][36] = 1;	doodle_right_transparency_texture[1][37] = 1;	doodle_right_transparency_texture[1][38] = 1;	doodle_right_transparency_texture[1][39] = 1;	doodle_right_transparency_texture[1][40] = 1;	doodle_right_transparency_texture[1][41] = 1;	doodle_right_transparency_texture[1][42] = 1;	doodle_right_transparency_texture[1][43] = 1;	doodle_right_transparency_texture[1][44] = 1;	doodle_right_transparency_texture[1][45] = 1;	doodle_right_transparency_texture[1][46] = 1;	doodle_right_transparency_texture[1][47] = 1;	doodle_right_transparency_texture[1][48] = 1;	doodle_right_transparency_texture[1][49] = 1;	doodle_right_transparency_texture[1][50] = 1;	doodle_right_transparency_texture[1][51] = 1;	doodle_right_transparency_texture[1][52] = 1;	doodle_right_transparency_texture[1][53] = 1;	doodle_right_transparency_texture[1][54] = 1;	doodle_right_transparency_texture[1][55] = 1;	doodle_right_transparency_texture[1][56] = 1;	doodle_right_transparency_texture[1][57] = 1;	doodle_right_transparency_texture[1][58] = 1;	doodle_right_transparency_texture[1][59] = 1;	doodle_right_transparency_texture[1][60] = 1;	doodle_right_transparency_texture[1][61] = 1;	doodle_right_transparency_texture[1][62] = 1;	doodle_right_transparency_texture[1][63] = 1;	doodle_right_transparency_texture[1][64] = 1;	doodle_right_transparency_texture[1][65] = 1;	doodle_right_transparency_texture[1][66] = 1;	doodle_right_transparency_texture[1][67] = 1;	doodle_right_transparency_texture[1][68] = 1;	doodle_right_transparency_texture[1][69] = 1;	doodle_right_transparency_texture[1][70] = 1;	doodle_right_transparency_texture[1][71] = 1;	doodle_right_transparency_texture[1][72] = 1;	doodle_right_transparency_texture[1][73] = 1;	doodle_right_transparency_texture[1][74] = 1;	doodle_right_transparency_texture[1][75] = 1;	doodle_right_transparency_texture[1][76] = 1;	doodle_right_transparency_texture[1][77] = 1;	doodle_right_transparency_texture[1][78] = 1;	doodle_right_transparency_texture[1][79] = 1;	doodle_right_transparency_texture[2][0] = 1;	doodle_right_transparency_texture[2][1] = 1;	doodle_right_transparency_texture[2][2] = 1;	doodle_right_transparency_texture[2][3] = 1;	doodle_right_transparency_texture[2][4] = 1;	doodle_right_transparency_texture[2][5] = 1;	doodle_right_transparency_texture[2][6] = 1;	doodle_right_transparency_texture[2][7] = 1;	doodle_right_transparency_texture[2][8] = 1;	doodle_right_transparency_texture[2][9] = 1;	doodle_right_transparency_texture[2][10] = 1;	doodle_right_transparency_texture[2][11] = 1;	doodle_right_transparency_texture[2][12] = 1;	doodle_right_transparency_texture[2][13] = 1;	doodle_right_transparency_texture[2][14] = 1;	doodle_right_transparency_texture[2][15] = 1;	doodle_right_transparency_texture[2][16] = 1;	doodle_right_transparency_texture[2][17] = 1;	doodle_right_transparency_texture[2][18] = 1;	doodle_right_transparency_texture[2][19] = 1;	doodle_right_transparency_texture[2][20] = 1;	doodle_right_transparency_texture[2][21] = 1;	doodle_right_transparency_texture[2][22] = 1;	doodle_right_transparency_texture[2][23] = 1;	doodle_right_transparency_texture[2][24] = 1;	doodle_right_transparency_texture[2][25] = 1;	doodle_right_transparency_texture[2][26] = 1;	doodle_right_transparency_texture[2][27] = 1;	doodle_right_transparency_texture[2][28] = 1;	doodle_right_transparency_texture[2][29] = 1;	doodle_right_transparency_texture[2][30] = 1;	doodle_right_transparency_texture[2][31] = 1;	doodle_right_transparency_texture[2][32] = 1;	doodle_right_transparency_texture[2][33] = 1;	doodle_right_transparency_texture[2][34] = 1;	doodle_right_transparency_texture[2][35] = 1;	doodle_right_transparency_texture[2][36] = 1;	doodle_right_transparency_texture[2][37] = 1;	doodle_right_transparency_texture[2][38] = 1;	doodle_right_transparency_texture[2][39] = 1;	doodle_right_transparency_texture[2][40] = 1;	doodle_right_transparency_texture[2][41] = 1;	doodle_right_transparency_texture[2][42] = 1;	doodle_right_transparency_texture[2][43] = 1;	doodle_right_transparency_texture[2][44] = 1;	doodle_right_transparency_texture[2][45] = 1;	doodle_right_transparency_texture[2][46] = 1;	doodle_right_transparency_texture[2][47] = 1;	doodle_right_transparency_texture[2][48] = 1;	doodle_right_transparency_texture[2][49] = 1;	doodle_right_transparency_texture[2][50] = 1;	doodle_right_transparency_texture[2][51] = 1;	doodle_right_transparency_texture[2][52] = 1;	doodle_right_transparency_texture[2][53] = 1;	doodle_right_transparency_texture[2][54] = 1;	doodle_right_transparency_texture[2][55] = 1;	doodle_right_transparency_texture[2][56] = 1;	doodle_right_transparency_texture[2][57] = 1;	doodle_right_transparency_texture[2][58] = 1;	doodle_right_transparency_texture[2][59] = 1;	doodle_right_transparency_texture[2][60] = 1;	doodle_right_transparency_texture[2][61] = 1;	doodle_right_transparency_texture[2][62] = 1;	doodle_right_transparency_texture[2][63] = 1;	doodle_right_transparency_texture[2][64] = 1;	doodle_right_transparency_texture[2][65] = 1;	doodle_right_transparency_texture[2][66] = 1;	doodle_right_transparency_texture[2][67] = 1;	doodle_right_transparency_texture[2][68] = 1;	doodle_right_transparency_texture[2][69] = 1;	doodle_right_transparency_texture[2][70] = 1;	doodle_right_transparency_texture[2][71] = 1;	doodle_right_transparency_texture[2][72] = 1;	doodle_right_transparency_texture[2][73] = 1;	doodle_right_transparency_texture[2][74] = 1;	doodle_right_transparency_texture[2][75] = 1;	doodle_right_transparency_texture[2][76] = 1;	doodle_right_transparency_texture[2][77] = 1;	doodle_right_transparency_texture[2][78] = 1;	doodle_right_transparency_texture[2][79] = 1;	doodle_right_transparency_texture[3][0] = 1;	doodle_right_transparency_texture[3][1] = 1;	doodle_right_transparency_texture[3][2] = 1;	doodle_right_transparency_texture[3][3] = 1;	doodle_right_transparency_texture[3][4] = 1;	doodle_right_transparency_texture[3][5] = 1;	doodle_right_transparency_texture[3][6] = 1;	doodle_right_transparency_texture[3][7] = 1;	doodle_right_transparency_texture[3][8] = 1;	doodle_right_transparency_texture[3][9] = 1;	doodle_right_transparency_texture[3][10] = 1;	doodle_right_transparency_texture[3][11] = 1;	doodle_right_transparency_texture[3][12] = 1;	doodle_right_transparency_texture[3][13] = 1;	doodle_right_transparency_texture[3][14] = 1;	doodle_right_transparency_texture[3][15] = 1;	doodle_right_transparency_texture[3][16] = 1;	doodle_right_transparency_texture[3][17] = 1;	doodle_right_transparency_texture[3][18] = 1;	doodle_right_transparency_texture[3][19] = 1;	doodle_right_transparency_texture[3][20] = 1;	doodle_right_transparency_texture[3][21] = 1;	doodle_right_transparency_texture[3][22] = 1;	doodle_right_transparency_texture[3][23] = 1;	doodle_right_transparency_texture[3][24] = 1;	doodle_right_transparency_texture[3][25] = 1;	doodle_right_transparency_texture[3][26] = 1;	doodle_right_transparency_texture[3][27] = 1;	doodle_right_transparency_texture[3][28] = 1;	doodle_right_transparency_texture[3][29] = 1;	doodle_right_transparency_texture[3][30] = 1;	doodle_right_transparency_texture[3][31] = 1;	doodle_right_transparency_texture[3][32] = 1;	doodle_right_transparency_texture[3][33] = 1;	doodle_right_transparency_texture[3][34] = 1;	doodle_right_transparency_texture[3][35] = 1;	doodle_right_transparency_texture[3][36] = 1;	doodle_right_transparency_texture[3][37] = 1;	doodle_right_transparency_texture[3][38] = 1;	doodle_right_transparency_texture[3][39] = 1;	doodle_right_transparency_texture[3][40] = 1;	doodle_right_transparency_texture[3][41] = 1;	doodle_right_transparency_texture[3][42] = 1;	doodle_right_transparency_texture[3][43] = 1;	doodle_right_transparency_texture[3][44] = 1;	doodle_right_transparency_texture[3][45] = 1;	doodle_right_transparency_texture[3][46] = 1;	doodle_right_transparency_texture[3][47] = 1;	doodle_right_transparency_texture[3][48] = 1;	doodle_right_transparency_texture[3][49] = 1;	doodle_right_transparency_texture[3][50] = 1;	doodle_right_transparency_texture[3][51] = 1;	doodle_right_transparency_texture[3][52] = 1;	doodle_right_transparency_texture[3][53] = 1;	doodle_right_transparency_texture[3][54] = 1;	doodle_right_transparency_texture[3][55] = 1;	doodle_right_transparency_texture[3][56] = 1;	doodle_right_transparency_texture[3][57] = 1;	doodle_right_transparency_texture[3][58] = 1;	doodle_right_transparency_texture[3][59] = 1;	doodle_right_transparency_texture[3][60] = 1;	doodle_right_transparency_texture[3][61] = 1;	doodle_right_transparency_texture[3][62] = 1;	doodle_right_transparency_texture[3][63] = 1;	doodle_right_transparency_texture[3][64] = 1;	doodle_right_transparency_texture[3][65] = 1;	doodle_right_transparency_texture[3][66] = 1;	doodle_right_transparency_texture[3][67] = 1;	doodle_right_transparency_texture[3][68] = 1;	doodle_right_transparency_texture[3][69] = 1;	doodle_right_transparency_texture[3][70] = 1;	doodle_right_transparency_texture[3][71] = 1;	doodle_right_transparency_texture[3][72] = 1;	doodle_right_transparency_texture[3][73] = 1;	doodle_right_transparency_texture[3][74] = 1;	doodle_right_transparency_texture[3][75] = 1;	doodle_right_transparency_texture[3][76] = 1;	doodle_right_transparency_texture[3][77] = 1;	doodle_right_transparency_texture[3][78] = 1;	doodle_right_transparency_texture[3][79] = 1;	doodle_right_transparency_texture[4][0] = 1;	doodle_right_transparency_texture[4][1] = 1;	doodle_right_transparency_texture[4][2] = 1;	doodle_right_transparency_texture[4][3] = 1;	doodle_right_transparency_texture[4][4] = 1;	doodle_right_transparency_texture[4][5] = 1;	doodle_right_transparency_texture[4][6] = 1;	doodle_right_transparency_texture[4][7] = 1;	doodle_right_transparency_texture[4][8] = 1;	doodle_right_transparency_texture[4][9] = 1;	doodle_right_transparency_texture[4][10] = 1;	doodle_right_transparency_texture[4][11] = 1;	doodle_right_transparency_texture[4][12] = 1;	doodle_right_transparency_texture[4][13] = 1;	doodle_right_transparency_texture[4][14] = 1;	doodle_right_transparency_texture[4][15] = 1;	doodle_right_transparency_texture[4][16] = 1;	doodle_right_transparency_texture[4][17] = 1;	doodle_right_transparency_texture[4][18] = 1;	doodle_right_transparency_texture[4][19] = 1;	doodle_right_transparency_texture[4][20] = 1;	doodle_right_transparency_texture[4][21] = 1;	doodle_right_transparency_texture[4][22] = 1;	doodle_right_transparency_texture[4][23] = 1;	doodle_right_transparency_texture[4][24] = 1;	doodle_right_transparency_texture[4][25] = 1;	doodle_right_transparency_texture[4][26] = 1;	doodle_right_transparency_texture[4][27] = 1;	doodle_right_transparency_texture[4][28] = 1;	doodle_right_transparency_texture[4][29] = 1;	doodle_right_transparency_texture[4][30] = 1;	doodle_right_transparency_texture[4][31] = 1;	doodle_right_transparency_texture[4][32] = 1;	doodle_right_transparency_texture[4][33] = 1;	doodle_right_transparency_texture[4][34] = 1;	doodle_right_transparency_texture[4][35] = 1;	doodle_right_transparency_texture[4][36] = 1;	doodle_right_transparency_texture[4][37] = 1;	doodle_right_transparency_texture[4][38] = 1;	doodle_right_transparency_texture[4][39] = 1;	doodle_right_transparency_texture[4][40] = 1;	doodle_right_transparency_texture[4][41] = 1;	doodle_right_transparency_texture[4][42] = 1;	doodle_right_transparency_texture[4][43] = 1;	doodle_right_transparency_texture[4][44] = 1;	doodle_right_transparency_texture[4][45] = 1;	doodle_right_transparency_texture[4][46] = 1;	doodle_right_transparency_texture[4][47] = 1;	doodle_right_transparency_texture[4][48] = 1;	doodle_right_transparency_texture[4][49] = 1;	doodle_right_transparency_texture[4][50] = 1;	doodle_right_transparency_texture[4][51] = 1;	doodle_right_transparency_texture[4][52] = 1;	doodle_right_transparency_texture[4][53] = 1;	doodle_right_transparency_texture[4][54] = 1;	doodle_right_transparency_texture[4][55] = 1;	doodle_right_transparency_texture[4][56] = 1;	doodle_right_transparency_texture[4][57] = 1;	doodle_right_transparency_texture[4][58] = 1;	doodle_right_transparency_texture[4][59] = 1;	doodle_right_transparency_texture[4][60] = 1;	doodle_right_transparency_texture[4][61] = 1;	doodle_right_transparency_texture[4][62] = 1;	doodle_right_transparency_texture[4][63] = 1;	doodle_right_transparency_texture[4][64] = 1;	doodle_right_transparency_texture[4][65] = 1;	doodle_right_transparency_texture[4][66] = 1;	doodle_right_transparency_texture[4][67] = 1;	doodle_right_transparency_texture[4][68] = 1;	doodle_right_transparency_texture[4][69] = 1;	doodle_right_transparency_texture[4][70] = 1;	doodle_right_transparency_texture[4][71] = 1;	doodle_right_transparency_texture[4][72] = 1;	doodle_right_transparency_texture[4][73] = 1;	doodle_right_transparency_texture[4][74] = 1;	doodle_right_transparency_texture[4][75] = 1;	doodle_right_transparency_texture[4][76] = 1;	doodle_right_transparency_texture[4][77] = 1;	doodle_right_transparency_texture[4][78] = 1;	doodle_right_transparency_texture[4][79] = 1;	doodle_right_transparency_texture[5][0] = 1;	doodle_right_transparency_texture[5][1] = 1;	doodle_right_transparency_texture[5][2] = 1;	doodle_right_transparency_texture[5][3] = 1;	doodle_right_transparency_texture[5][4] = 1;	doodle_right_transparency_texture[5][5] = 1;	doodle_right_transparency_texture[5][6] = 1;	doodle_right_transparency_texture[5][7] = 1;	doodle_right_transparency_texture[5][8] = 1;	doodle_right_transparency_texture[5][9] = 1;	doodle_right_transparency_texture[5][10] = 1;	doodle_right_transparency_texture[5][11] = 1;	doodle_right_transparency_texture[5][12] = 1;	doodle_right_transparency_texture[5][13] = 1;	doodle_right_transparency_texture[5][14] = 1;	doodle_right_transparency_texture[5][15] = 1;	doodle_right_transparency_texture[5][16] = 1;	doodle_right_transparency_texture[5][17] = 1;	doodle_right_transparency_texture[5][18] = 1;	doodle_right_transparency_texture[5][19] = 1;	doodle_right_transparency_texture[5][20] = 1;	doodle_right_transparency_texture[5][21] = 1;	doodle_right_transparency_texture[5][22] = 1;	doodle_right_transparency_texture[5][23] = 1;	doodle_right_transparency_texture[5][24] = 1;	doodle_right_transparency_texture[5][25] = 1;	doodle_right_transparency_texture[5][26] = 1;	doodle_right_transparency_texture[5][27] = 1;	doodle_right_transparency_texture[5][28] = 1;	doodle_right_transparency_texture[5][29] = 1;	doodle_right_transparency_texture[5][30] = 1;	doodle_right_transparency_texture[5][31] = 1;	doodle_right_transparency_texture[5][32] = 1;	doodle_right_transparency_texture[5][33] = 1;	doodle_right_transparency_texture[5][34] = 1;	doodle_right_transparency_texture[5][35] = 1;	doodle_right_transparency_texture[5][36] = 1;	doodle_right_transparency_texture[5][37] = 1;	doodle_right_transparency_texture[5][38] = 1;	doodle_right_transparency_texture[5][39] = 1;	doodle_right_transparency_texture[5][40] = 1;	doodle_right_transparency_texture[5][41] = 1;	doodle_right_transparency_texture[5][42] = 1;	doodle_right_transparency_texture[5][43] = 1;	doodle_right_transparency_texture[5][44] = 1;	doodle_right_transparency_texture[5][45] = 1;	doodle_right_transparency_texture[5][46] = 1;	doodle_right_transparency_texture[5][47] = 1;	doodle_right_transparency_texture[5][48] = 1;	doodle_right_transparency_texture[5][49] = 1;	doodle_right_transparency_texture[5][50] = 1;	doodle_right_transparency_texture[5][51] = 1;	doodle_right_transparency_texture[5][52] = 1;	doodle_right_transparency_texture[5][53] = 1;	doodle_right_transparency_texture[5][54] = 1;	doodle_right_transparency_texture[5][55] = 1;	doodle_right_transparency_texture[5][56] = 1;	doodle_right_transparency_texture[5][57] = 1;	doodle_right_transparency_texture[5][58] = 1;	doodle_right_transparency_texture[5][59] = 1;	doodle_right_transparency_texture[5][60] = 1;	doodle_right_transparency_texture[5][61] = 1;	doodle_right_transparency_texture[5][62] = 1;	doodle_right_transparency_texture[5][63] = 1;	doodle_right_transparency_texture[5][64] = 1;	doodle_right_transparency_texture[5][65] = 1;	doodle_right_transparency_texture[5][66] = 1;	doodle_right_transparency_texture[5][67] = 1;	doodle_right_transparency_texture[5][68] = 1;	doodle_right_transparency_texture[5][69] = 1;	doodle_right_transparency_texture[5][70] = 1;	doodle_right_transparency_texture[5][71] = 1;	doodle_right_transparency_texture[5][72] = 1;	doodle_right_transparency_texture[5][73] = 1;	doodle_right_transparency_texture[5][74] = 1;	doodle_right_transparency_texture[5][75] = 1;	doodle_right_transparency_texture[5][76] = 1;	doodle_right_transparency_texture[5][77] = 1;	doodle_right_transparency_texture[5][78] = 1;	doodle_right_transparency_texture[5][79] = 1;	doodle_right_transparency_texture[6][0] = 1;	doodle_right_transparency_texture[6][1] = 1;	doodle_right_transparency_texture[6][2] = 1;	doodle_right_transparency_texture[6][3] = 1;	doodle_right_transparency_texture[6][4] = 1;	doodle_right_transparency_texture[6][5] = 1;	doodle_right_transparency_texture[6][6] = 1;	doodle_right_transparency_texture[6][7] = 1;	doodle_right_transparency_texture[6][8] = 1;	doodle_right_transparency_texture[6][9] = 1;	doodle_right_transparency_texture[6][10] = 1;	doodle_right_transparency_texture[6][11] = 1;	doodle_right_transparency_texture[6][12] = 1;	doodle_right_transparency_texture[6][13] = 1;	doodle_right_transparency_texture[6][14] = 1;	doodle_right_transparency_texture[6][15] = 1;	doodle_right_transparency_texture[6][16] = 1;	doodle_right_transparency_texture[6][17] = 1;	doodle_right_transparency_texture[6][18] = 1;	doodle_right_transparency_texture[6][19] = 1;	doodle_right_transparency_texture[6][20] = 1;	doodle_right_transparency_texture[6][21] = 1;	doodle_right_transparency_texture[6][22] = 1;	doodle_right_transparency_texture[6][23] = 1;	doodle_right_transparency_texture[6][24] = 1;	doodle_right_transparency_texture[6][25] = 1;	doodle_right_transparency_texture[6][26] = 1;	doodle_right_transparency_texture[6][27] = 1;	doodle_right_transparency_texture[6][28] = 1;	doodle_right_transparency_texture[6][29] = 1;	doodle_right_transparency_texture[6][30] = 1;	doodle_right_transparency_texture[6][31] = 1;	doodle_right_transparency_texture[6][32] = 1;	doodle_right_transparency_texture[6][33] = 1;	doodle_right_transparency_texture[6][34] = 1;	doodle_right_transparency_texture[6][35] = 1;	doodle_right_transparency_texture[6][36] = 1;	doodle_right_transparency_texture[6][37] = 1;	doodle_right_transparency_texture[6][38] = 1;	doodle_right_transparency_texture[6][39] = 1;	doodle_right_transparency_texture[6][40] = 1;	doodle_right_transparency_texture[6][41] = 1;	doodle_right_transparency_texture[6][42] = 1;	doodle_right_transparency_texture[6][43] = 1;	doodle_right_transparency_texture[6][44] = 1;	doodle_right_transparency_texture[6][45] = 1;	doodle_right_transparency_texture[6][46] = 1;	doodle_right_transparency_texture[6][47] = 1;	doodle_right_transparency_texture[6][48] = 1;	doodle_right_transparency_texture[6][49] = 1;	doodle_right_transparency_texture[6][50] = 1;	doodle_right_transparency_texture[6][51] = 1;	doodle_right_transparency_texture[6][52] = 1;	doodle_right_transparency_texture[6][53] = 1;	doodle_right_transparency_texture[6][54] = 1;	doodle_right_transparency_texture[6][55] = 1;	doodle_right_transparency_texture[6][56] = 1;	doodle_right_transparency_texture[6][57] = 1;	doodle_right_transparency_texture[6][58] = 1;	doodle_right_transparency_texture[6][59] = 1;	doodle_right_transparency_texture[6][60] = 1;	doodle_right_transparency_texture[6][61] = 1;	doodle_right_transparency_texture[6][62] = 1;	doodle_right_transparency_texture[6][63] = 1;	doodle_right_transparency_texture[6][64] = 1;	doodle_right_transparency_texture[6][65] = 1;	doodle_right_transparency_texture[6][66] = 1;	doodle_right_transparency_texture[6][67] = 1;	doodle_right_transparency_texture[6][68] = 1;	doodle_right_transparency_texture[6][69] = 1;	doodle_right_transparency_texture[6][70] = 1;	doodle_right_transparency_texture[6][71] = 1;	doodle_right_transparency_texture[6][72] = 1;	doodle_right_transparency_texture[6][73] = 1;	doodle_right_transparency_texture[6][74] = 1;	doodle_right_transparency_texture[6][75] = 1;	doodle_right_transparency_texture[6][76] = 1;	doodle_right_transparency_texture[6][77] = 1;	doodle_right_transparency_texture[6][78] = 1;	doodle_right_transparency_texture[6][79] = 1;	doodle_right_transparency_texture[7][0] = 1;	doodle_right_transparency_texture[7][1] = 1;	doodle_right_transparency_texture[7][2] = 1;	doodle_right_transparency_texture[7][3] = 1;	doodle_right_transparency_texture[7][4] = 1;	doodle_right_transparency_texture[7][5] = 1;	doodle_right_transparency_texture[7][6] = 1;	doodle_right_transparency_texture[7][7] = 1;	doodle_right_transparency_texture[7][8] = 1;	doodle_right_transparency_texture[7][9] = 1;	doodle_right_transparency_texture[7][10] = 1;	doodle_right_transparency_texture[7][11] = 1;	doodle_right_transparency_texture[7][12] = 1;	doodle_right_transparency_texture[7][13] = 1;	doodle_right_transparency_texture[7][14] = 1;	doodle_right_transparency_texture[7][15] = 1;	doodle_right_transparency_texture[7][16] = 1;	doodle_right_transparency_texture[7][17] = 1;	doodle_right_transparency_texture[7][18] = 1;	doodle_right_transparency_texture[7][19] = 1;	doodle_right_transparency_texture[7][20] = 1;	doodle_right_transparency_texture[7][21] = 1;	doodle_right_transparency_texture[7][22] = 1;	doodle_right_transparency_texture[7][23] = 1;	doodle_right_transparency_texture[7][24] = 1;	doodle_right_transparency_texture[7][25] = 1;	doodle_right_transparency_texture[7][26] = 1;	doodle_right_transparency_texture[7][27] = 1;	doodle_right_transparency_texture[7][28] = 1;	doodle_right_transparency_texture[7][29] = 1;	doodle_right_transparency_texture[7][30] = 1;	doodle_right_transparency_texture[7][31] = 1;	doodle_right_transparency_texture[7][32] = 1;	doodle_right_transparency_texture[7][33] = 1;	doodle_right_transparency_texture[7][34] = 1;	doodle_right_transparency_texture[7][35] = 1;	doodle_right_transparency_texture[7][36] = 1;	doodle_right_transparency_texture[7][37] = 1;	doodle_right_transparency_texture[7][38] = 1;	doodle_right_transparency_texture[7][39] = 1;	doodle_right_transparency_texture[7][40] = 1;	doodle_right_transparency_texture[7][41] = 1;	doodle_right_transparency_texture[7][42] = 1;	doodle_right_transparency_texture[7][43] = 1;	doodle_right_transparency_texture[7][44] = 1;	doodle_right_transparency_texture[7][45] = 1;	doodle_right_transparency_texture[7][46] = 1;	doodle_right_transparency_texture[7][47] = 1;	doodle_right_transparency_texture[7][48] = 1;	doodle_right_transparency_texture[7][49] = 1;	doodle_right_transparency_texture[7][50] = 1;	doodle_right_transparency_texture[7][51] = 1;	doodle_right_transparency_texture[7][52] = 1;	doodle_right_transparency_texture[7][53] = 1;	doodle_right_transparency_texture[7][54] = 1;	doodle_right_transparency_texture[7][55] = 1;	doodle_right_transparency_texture[7][56] = 1;	doodle_right_transparency_texture[7][57] = 1;	doodle_right_transparency_texture[7][58] = 1;	doodle_right_transparency_texture[7][59] = 1;	doodle_right_transparency_texture[7][60] = 1;	doodle_right_transparency_texture[7][61] = 1;	doodle_right_transparency_texture[7][62] = 1;	doodle_right_transparency_texture[7][63] = 1;	doodle_right_transparency_texture[7][64] = 1;	doodle_right_transparency_texture[7][65] = 1;	doodle_right_transparency_texture[7][66] = 1;	doodle_right_transparency_texture[7][67] = 1;	doodle_right_transparency_texture[7][68] = 1;	doodle_right_transparency_texture[7][69] = 1;	doodle_right_transparency_texture[7][70] = 1;	doodle_right_transparency_texture[7][71] = 1;	doodle_right_transparency_texture[7][72] = 1;	doodle_right_transparency_texture[7][73] = 1;	doodle_right_transparency_texture[7][74] = 1;	doodle_right_transparency_texture[7][75] = 1;	doodle_right_transparency_texture[7][76] = 1;	doodle_right_transparency_texture[7][77] = 1;	doodle_right_transparency_texture[7][78] = 1;	doodle_right_transparency_texture[7][79] = 1;	doodle_right_transparency_texture[8][0] = 1;	doodle_right_transparency_texture[8][1] = 1;	doodle_right_transparency_texture[8][2] = 1;	doodle_right_transparency_texture[8][3] = 1;	doodle_right_transparency_texture[8][4] = 1;	doodle_right_transparency_texture[8][5] = 1;	doodle_right_transparency_texture[8][6] = 1;	doodle_right_transparency_texture[8][7] = 1;	doodle_right_transparency_texture[8][8] = 1;	doodle_right_transparency_texture[8][9] = 1;	doodle_right_transparency_texture[8][10] = 1;	doodle_right_transparency_texture[8][11] = 1;	doodle_right_transparency_texture[8][12] = 0;	doodle_right_transparency_texture[8][13] = 0;	doodle_right_transparency_texture[8][14] = 0;	doodle_right_transparency_texture[8][15] = 0;	doodle_right_transparency_texture[8][16] = 0;	doodle_right_transparency_texture[8][17] = 0;	doodle_right_transparency_texture[8][18] = 0;	doodle_right_transparency_texture[8][19] = 0;	doodle_right_transparency_texture[8][20] = 0;	doodle_right_transparency_texture[8][21] = 0;	doodle_right_transparency_texture[8][22] = 0;	doodle_right_transparency_texture[8][23] = 0;	doodle_right_transparency_texture[8][24] = 0;	doodle_right_transparency_texture[8][25] = 0;	doodle_right_transparency_texture[8][26] = 0;	doodle_right_transparency_texture[8][27] = 0;	doodle_right_transparency_texture[8][28] = 0;	doodle_right_transparency_texture[8][29] = 0;	doodle_right_transparency_texture[8][30] = 0;	doodle_right_transparency_texture[8][31] = 0;	doodle_right_transparency_texture[8][32] = 0;	doodle_right_transparency_texture[8][33] = 0;	doodle_right_transparency_texture[8][34] = 0;	doodle_right_transparency_texture[8][35] = 0;	doodle_right_transparency_texture[8][36] = 0;	doodle_right_transparency_texture[8][37] = 0;	doodle_right_transparency_texture[8][38] = 0;	doodle_right_transparency_texture[8][39] = 0;	doodle_right_transparency_texture[8][40] = 0;	doodle_right_transparency_texture[8][41] = 0;	doodle_right_transparency_texture[8][42] = 0;	doodle_right_transparency_texture[8][43] = 0;	doodle_right_transparency_texture[8][44] = 1;	doodle_right_transparency_texture[8][45] = 1;	doodle_right_transparency_texture[8][46] = 1;	doodle_right_transparency_texture[8][47] = 1;	doodle_right_transparency_texture[8][48] = 1;	doodle_right_transparency_texture[8][49] = 1;	doodle_right_transparency_texture[8][50] = 1;	doodle_right_transparency_texture[8][51] = 1;	doodle_right_transparency_texture[8][52] = 1;	doodle_right_transparency_texture[8][53] = 1;	doodle_right_transparency_texture[8][54] = 1;	doodle_right_transparency_texture[8][55] = 1;	doodle_right_transparency_texture[8][56] = 1;	doodle_right_transparency_texture[8][57] = 1;	doodle_right_transparency_texture[8][58] = 1;	doodle_right_transparency_texture[8][59] = 1;	doodle_right_transparency_texture[8][60] = 1;	doodle_right_transparency_texture[8][61] = 1;	doodle_right_transparency_texture[8][62] = 1;	doodle_right_transparency_texture[8][63] = 1;	doodle_right_transparency_texture[8][64] = 1;	doodle_right_transparency_texture[8][65] = 1;	doodle_right_transparency_texture[8][66] = 1;	doodle_right_transparency_texture[8][67] = 1;	doodle_right_transparency_texture[8][68] = 1;	doodle_right_transparency_texture[8][69] = 1;	doodle_right_transparency_texture[8][70] = 1;	doodle_right_transparency_texture[8][71] = 1;	doodle_right_transparency_texture[8][72] = 1;	doodle_right_transparency_texture[8][73] = 1;	doodle_right_transparency_texture[8][74] = 1;	doodle_right_transparency_texture[8][75] = 1;	doodle_right_transparency_texture[8][76] = 1;	doodle_right_transparency_texture[8][77] = 1;	doodle_right_transparency_texture[8][78] = 1;	doodle_right_transparency_texture[8][79] = 1;	doodle_right_transparency_texture[9][0] = 1;	doodle_right_transparency_texture[9][1] = 1;	doodle_right_transparency_texture[9][2] = 1;	doodle_right_transparency_texture[9][3] = 1;	doodle_right_transparency_texture[9][4] = 1;	doodle_right_transparency_texture[9][5] = 1;	doodle_right_transparency_texture[9][6] = 1;	doodle_right_transparency_texture[9][7] = 1;	doodle_right_transparency_texture[9][8] = 1;	doodle_right_transparency_texture[9][9] = 1;	doodle_right_transparency_texture[9][10] = 1;	doodle_right_transparency_texture[9][11] = 1;	doodle_right_transparency_texture[9][12] = 0;	doodle_right_transparency_texture[9][13] = 0;	doodle_right_transparency_texture[9][14] = 0;	doodle_right_transparency_texture[9][15] = 0;	doodle_right_transparency_texture[9][16] = 0;	doodle_right_transparency_texture[9][17] = 0;	doodle_right_transparency_texture[9][18] = 0;	doodle_right_transparency_texture[9][19] = 0;	doodle_right_transparency_texture[9][20] = 0;	doodle_right_transparency_texture[9][21] = 0;	doodle_right_transparency_texture[9][22] = 0;	doodle_right_transparency_texture[9][23] = 0;	doodle_right_transparency_texture[9][24] = 0;	doodle_right_transparency_texture[9][25] = 0;	doodle_right_transparency_texture[9][26] = 0;	doodle_right_transparency_texture[9][27] = 0;	doodle_right_transparency_texture[9][28] = 0;	doodle_right_transparency_texture[9][29] = 0;	doodle_right_transparency_texture[9][30] = 0;	doodle_right_transparency_texture[9][31] = 0;	doodle_right_transparency_texture[9][32] = 0;	doodle_right_transparency_texture[9][33] = 0;	doodle_right_transparency_texture[9][34] = 0;	doodle_right_transparency_texture[9][35] = 0;	doodle_right_transparency_texture[9][36] = 0;	doodle_right_transparency_texture[9][37] = 0;	doodle_right_transparency_texture[9][38] = 0;	doodle_right_transparency_texture[9][39] = 0;	doodle_right_transparency_texture[9][40] = 0;	doodle_right_transparency_texture[9][41] = 0;	doodle_right_transparency_texture[9][42] = 0;	doodle_right_transparency_texture[9][43] = 0;	doodle_right_transparency_texture[9][44] = 1;	doodle_right_transparency_texture[9][45] = 1;	doodle_right_transparency_texture[9][46] = 1;	doodle_right_transparency_texture[9][47] = 1;	doodle_right_transparency_texture[9][48] = 1;	doodle_right_transparency_texture[9][49] = 1;	doodle_right_transparency_texture[9][50] = 1;	doodle_right_transparency_texture[9][51] = 1;	doodle_right_transparency_texture[9][52] = 1;	doodle_right_transparency_texture[9][53] = 1;	doodle_right_transparency_texture[9][54] = 1;	doodle_right_transparency_texture[9][55] = 1;	doodle_right_transparency_texture[9][56] = 1;	doodle_right_transparency_texture[9][57] = 1;	doodle_right_transparency_texture[9][58] = 1;	doodle_right_transparency_texture[9][59] = 1;	doodle_right_transparency_texture[9][60] = 1;	doodle_right_transparency_texture[9][61] = 1;	doodle_right_transparency_texture[9][62] = 1;	doodle_right_transparency_texture[9][63] = 1;	doodle_right_transparency_texture[9][64] = 1;	doodle_right_transparency_texture[9][65] = 1;	doodle_right_transparency_texture[9][66] = 1;	doodle_right_transparency_texture[9][67] = 1;	doodle_right_transparency_texture[9][68] = 1;	doodle_right_transparency_texture[9][69] = 1;	doodle_right_transparency_texture[9][70] = 1;	doodle_right_transparency_texture[9][71] = 1;	doodle_right_transparency_texture[9][72] = 1;	doodle_right_transparency_texture[9][73] = 1;	doodle_right_transparency_texture[9][74] = 1;	doodle_right_transparency_texture[9][75] = 1;	doodle_right_transparency_texture[9][76] = 1;	doodle_right_transparency_texture[9][77] = 1;	doodle_right_transparency_texture[9][78] = 1;	doodle_right_transparency_texture[9][79] = 1;	doodle_right_transparency_texture[10][0] = 1;	doodle_right_transparency_texture[10][1] = 1;	doodle_right_transparency_texture[10][2] = 1;	doodle_right_transparency_texture[10][3] = 1;	doodle_right_transparency_texture[10][4] = 1;	doodle_right_transparency_texture[10][5] = 1;	doodle_right_transparency_texture[10][6] = 1;	doodle_right_transparency_texture[10][7] = 1;	doodle_right_transparency_texture[10][8] = 1;	doodle_right_transparency_texture[10][9] = 1;	doodle_right_transparency_texture[10][10] = 1;	doodle_right_transparency_texture[10][11] = 1;	doodle_right_transparency_texture[10][12] = 0;	doodle_right_transparency_texture[10][13] = 0;	doodle_right_transparency_texture[10][14] = 0;	doodle_right_transparency_texture[10][15] = 0;	doodle_right_transparency_texture[10][16] = 0;	doodle_right_transparency_texture[10][17] = 0;	doodle_right_transparency_texture[10][18] = 0;	doodle_right_transparency_texture[10][19] = 0;	doodle_right_transparency_texture[10][20] = 0;	doodle_right_transparency_texture[10][21] = 0;	doodle_right_transparency_texture[10][22] = 0;	doodle_right_transparency_texture[10][23] = 0;	doodle_right_transparency_texture[10][24] = 0;	doodle_right_transparency_texture[10][25] = 0;	doodle_right_transparency_texture[10][26] = 0;	doodle_right_transparency_texture[10][27] = 0;	doodle_right_transparency_texture[10][28] = 0;	doodle_right_transparency_texture[10][29] = 0;	doodle_right_transparency_texture[10][30] = 0;	doodle_right_transparency_texture[10][31] = 0;	doodle_right_transparency_texture[10][32] = 0;	doodle_right_transparency_texture[10][33] = 0;	doodle_right_transparency_texture[10][34] = 0;	doodle_right_transparency_texture[10][35] = 0;	doodle_right_transparency_texture[10][36] = 0;	doodle_right_transparency_texture[10][37] = 0;	doodle_right_transparency_texture[10][38] = 0;	doodle_right_transparency_texture[10][39] = 0;	doodle_right_transparency_texture[10][40] = 0;	doodle_right_transparency_texture[10][41] = 0;	doodle_right_transparency_texture[10][42] = 0;	doodle_right_transparency_texture[10][43] = 0;	doodle_right_transparency_texture[10][44] = 1;	doodle_right_transparency_texture[10][45] = 1;	doodle_right_transparency_texture[10][46] = 1;	doodle_right_transparency_texture[10][47] = 1;	doodle_right_transparency_texture[10][48] = 1;	doodle_right_transparency_texture[10][49] = 1;	doodle_right_transparency_texture[10][50] = 1;	doodle_right_transparency_texture[10][51] = 1;	doodle_right_transparency_texture[10][52] = 1;	doodle_right_transparency_texture[10][53] = 1;	doodle_right_transparency_texture[10][54] = 1;	doodle_right_transparency_texture[10][55] = 1;	doodle_right_transparency_texture[10][56] = 1;	doodle_right_transparency_texture[10][57] = 1;	doodle_right_transparency_texture[10][58] = 1;	doodle_right_transparency_texture[10][59] = 1;	doodle_right_transparency_texture[10][60] = 1;	doodle_right_transparency_texture[10][61] = 1;	doodle_right_transparency_texture[10][62] = 1;	doodle_right_transparency_texture[10][63] = 1;	doodle_right_transparency_texture[10][64] = 1;	doodle_right_transparency_texture[10][65] = 1;	doodle_right_transparency_texture[10][66] = 1;	doodle_right_transparency_texture[10][67] = 1;	doodle_right_transparency_texture[10][68] = 1;	doodle_right_transparency_texture[10][69] = 1;	doodle_right_transparency_texture[10][70] = 1;	doodle_right_transparency_texture[10][71] = 1;	doodle_right_transparency_texture[10][72] = 1;	doodle_right_transparency_texture[10][73] = 1;	doodle_right_transparency_texture[10][74] = 1;	doodle_right_transparency_texture[10][75] = 1;	doodle_right_transparency_texture[10][76] = 1;	doodle_right_transparency_texture[10][77] = 1;	doodle_right_transparency_texture[10][78] = 1;	doodle_right_transparency_texture[10][79] = 1;	doodle_right_transparency_texture[11][0] = 1;	doodle_right_transparency_texture[11][1] = 1;	doodle_right_transparency_texture[11][2] = 1;	doodle_right_transparency_texture[11][3] = 1;	doodle_right_transparency_texture[11][4] = 1;	doodle_right_transparency_texture[11][5] = 1;	doodle_right_transparency_texture[11][6] = 1;	doodle_right_transparency_texture[11][7] = 1;	doodle_right_transparency_texture[11][8] = 1;	doodle_right_transparency_texture[11][9] = 1;	doodle_right_transparency_texture[11][10] = 1;	doodle_right_transparency_texture[11][11] = 1;	doodle_right_transparency_texture[11][12] = 0;	doodle_right_transparency_texture[11][13] = 0;	doodle_right_transparency_texture[11][14] = 0;	doodle_right_transparency_texture[11][15] = 0;	doodle_right_transparency_texture[11][16] = 0;	doodle_right_transparency_texture[11][17] = 0;	doodle_right_transparency_texture[11][18] = 0;	doodle_right_transparency_texture[11][19] = 0;	doodle_right_transparency_texture[11][20] = 0;	doodle_right_transparency_texture[11][21] = 0;	doodle_right_transparency_texture[11][22] = 0;	doodle_right_transparency_texture[11][23] = 0;	doodle_right_transparency_texture[11][24] = 0;	doodle_right_transparency_texture[11][25] = 0;	doodle_right_transparency_texture[11][26] = 0;	doodle_right_transparency_texture[11][27] = 0;	doodle_right_transparency_texture[11][28] = 0;	doodle_right_transparency_texture[11][29] = 0;	doodle_right_transparency_texture[11][30] = 0;	doodle_right_transparency_texture[11][31] = 0;	doodle_right_transparency_texture[11][32] = 0;	doodle_right_transparency_texture[11][33] = 0;	doodle_right_transparency_texture[11][34] = 0;	doodle_right_transparency_texture[11][35] = 0;	doodle_right_transparency_texture[11][36] = 0;	doodle_right_transparency_texture[11][37] = 0;	doodle_right_transparency_texture[11][38] = 0;	doodle_right_transparency_texture[11][39] = 0;	doodle_right_transparency_texture[11][40] = 0;	doodle_right_transparency_texture[11][41] = 0;	doodle_right_transparency_texture[11][42] = 0;	doodle_right_transparency_texture[11][43] = 0;	doodle_right_transparency_texture[11][44] = 1;	doodle_right_transparency_texture[11][45] = 1;	doodle_right_transparency_texture[11][46] = 1;	doodle_right_transparency_texture[11][47] = 1;	doodle_right_transparency_texture[11][48] = 1;	doodle_right_transparency_texture[11][49] = 1;	doodle_right_transparency_texture[11][50] = 1;	doodle_right_transparency_texture[11][51] = 1;	doodle_right_transparency_texture[11][52] = 1;	doodle_right_transparency_texture[11][53] = 1;	doodle_right_transparency_texture[11][54] = 1;	doodle_right_transparency_texture[11][55] = 1;	doodle_right_transparency_texture[11][56] = 1;	doodle_right_transparency_texture[11][57] = 1;	doodle_right_transparency_texture[11][58] = 1;	doodle_right_transparency_texture[11][59] = 1;	doodle_right_transparency_texture[11][60] = 1;	doodle_right_transparency_texture[11][61] = 1;	doodle_right_transparency_texture[11][62] = 1;	doodle_right_transparency_texture[11][63] = 1;	doodle_right_transparency_texture[11][64] = 1;	doodle_right_transparency_texture[11][65] = 1;	doodle_right_transparency_texture[11][66] = 1;	doodle_right_transparency_texture[11][67] = 1;	doodle_right_transparency_texture[11][68] = 1;	doodle_right_transparency_texture[11][69] = 1;	doodle_right_transparency_texture[11][70] = 1;	doodle_right_transparency_texture[11][71] = 1;	doodle_right_transparency_texture[11][72] = 1;	doodle_right_transparency_texture[11][73] = 1;	doodle_right_transparency_texture[11][74] = 1;	doodle_right_transparency_texture[11][75] = 1;	doodle_right_transparency_texture[11][76] = 1;	doodle_right_transparency_texture[11][77] = 1;	doodle_right_transparency_texture[11][78] = 1;	doodle_right_transparency_texture[11][79] = 1;	doodle_right_transparency_texture[12][0] = 1;	doodle_right_transparency_texture[12][1] = 1;	doodle_right_transparency_texture[12][2] = 1;	doodle_right_transparency_texture[12][3] = 1;	doodle_right_transparency_texture[12][4] = 1;	doodle_right_transparency_texture[12][5] = 1;	doodle_right_transparency_texture[12][6] = 1;	doodle_right_transparency_texture[12][7] = 1;	doodle_right_transparency_texture[12][8] = 0;	doodle_right_transparency_texture[12][9] = 0;	doodle_right_transparency_texture[12][10] = 0;	doodle_right_transparency_texture[12][11] = 0;	doodle_right_transparency_texture[12][12] = 0;	doodle_right_transparency_texture[12][13] = 0;	doodle_right_transparency_texture[12][14] = 0;	doodle_right_transparency_texture[12][15] = 0;	doodle_right_transparency_texture[12][16] = 0;	doodle_right_transparency_texture[12][17] = 0;	doodle_right_transparency_texture[12][18] = 0;	doodle_right_transparency_texture[12][19] = 0;	doodle_right_transparency_texture[12][20] = 0;	doodle_right_transparency_texture[12][21] = 0;	doodle_right_transparency_texture[12][22] = 0;	doodle_right_transparency_texture[12][23] = 0;	doodle_right_transparency_texture[12][24] = 0;	doodle_right_transparency_texture[12][25] = 0;	doodle_right_transparency_texture[12][26] = 0;	doodle_right_transparency_texture[12][27] = 0;	doodle_right_transparency_texture[12][28] = 0;	doodle_right_transparency_texture[12][29] = 0;	doodle_right_transparency_texture[12][30] = 0;	doodle_right_transparency_texture[12][31] = 0;	doodle_right_transparency_texture[12][32] = 0;	doodle_right_transparency_texture[12][33] = 0;	doodle_right_transparency_texture[12][34] = 0;	doodle_right_transparency_texture[12][35] = 0;	doodle_right_transparency_texture[12][36] = 0;	doodle_right_transparency_texture[12][37] = 0;	doodle_right_transparency_texture[12][38] = 0;	doodle_right_transparency_texture[12][39] = 0;	doodle_right_transparency_texture[12][40] = 0;	doodle_right_transparency_texture[12][41] = 0;	doodle_right_transparency_texture[12][42] = 0;	doodle_right_transparency_texture[12][43] = 0;	doodle_right_transparency_texture[12][44] = 0;	doodle_right_transparency_texture[12][45] = 0;	doodle_right_transparency_texture[12][46] = 0;	doodle_right_transparency_texture[12][47] = 0;	doodle_right_transparency_texture[12][48] = 1;	doodle_right_transparency_texture[12][49] = 1;	doodle_right_transparency_texture[12][50] = 1;	doodle_right_transparency_texture[12][51] = 1;	doodle_right_transparency_texture[12][52] = 1;	doodle_right_transparency_texture[12][53] = 1;	doodle_right_transparency_texture[12][54] = 1;	doodle_right_transparency_texture[12][55] = 1;	doodle_right_transparency_texture[12][56] = 1;	doodle_right_transparency_texture[12][57] = 1;	doodle_right_transparency_texture[12][58] = 1;	doodle_right_transparency_texture[12][59] = 1;	doodle_right_transparency_texture[12][60] = 1;	doodle_right_transparency_texture[12][61] = 1;	doodle_right_transparency_texture[12][62] = 1;	doodle_right_transparency_texture[12][63] = 1;	doodle_right_transparency_texture[12][64] = 1;	doodle_right_transparency_texture[12][65] = 1;	doodle_right_transparency_texture[12][66] = 1;	doodle_right_transparency_texture[12][67] = 1;	doodle_right_transparency_texture[12][68] = 1;	doodle_right_transparency_texture[12][69] = 1;	doodle_right_transparency_texture[12][70] = 1;	doodle_right_transparency_texture[12][71] = 1;	doodle_right_transparency_texture[12][72] = 1;	doodle_right_transparency_texture[12][73] = 1;	doodle_right_transparency_texture[12][74] = 1;	doodle_right_transparency_texture[12][75] = 1;	doodle_right_transparency_texture[12][76] = 1;	doodle_right_transparency_texture[12][77] = 1;	doodle_right_transparency_texture[12][78] = 1;	doodle_right_transparency_texture[12][79] = 1;	doodle_right_transparency_texture[13][0] = 1;	doodle_right_transparency_texture[13][1] = 1;	doodle_right_transparency_texture[13][2] = 1;	doodle_right_transparency_texture[13][3] = 1;	doodle_right_transparency_texture[13][4] = 1;	doodle_right_transparency_texture[13][5] = 1;	doodle_right_transparency_texture[13][6] = 1;	doodle_right_transparency_texture[13][7] = 1;	doodle_right_transparency_texture[13][8] = 0;	doodle_right_transparency_texture[13][9] = 0;	doodle_right_transparency_texture[13][10] = 0;	doodle_right_transparency_texture[13][11] = 0;	doodle_right_transparency_texture[13][12] = 0;	doodle_right_transparency_texture[13][13] = 0;	doodle_right_transparency_texture[13][14] = 0;	doodle_right_transparency_texture[13][15] = 0;	doodle_right_transparency_texture[13][16] = 0;	doodle_right_transparency_texture[13][17] = 0;	doodle_right_transparency_texture[13][18] = 0;	doodle_right_transparency_texture[13][19] = 0;	doodle_right_transparency_texture[13][20] = 0;	doodle_right_transparency_texture[13][21] = 0;	doodle_right_transparency_texture[13][22] = 0;	doodle_right_transparency_texture[13][23] = 0;	doodle_right_transparency_texture[13][24] = 0;	doodle_right_transparency_texture[13][25] = 0;	doodle_right_transparency_texture[13][26] = 0;	doodle_right_transparency_texture[13][27] = 0;	doodle_right_transparency_texture[13][28] = 0;	doodle_right_transparency_texture[13][29] = 0;	doodle_right_transparency_texture[13][30] = 0;	doodle_right_transparency_texture[13][31] = 0;	doodle_right_transparency_texture[13][32] = 0;	doodle_right_transparency_texture[13][33] = 0;	doodle_right_transparency_texture[13][34] = 0;	doodle_right_transparency_texture[13][35] = 0;	doodle_right_transparency_texture[13][36] = 0;	doodle_right_transparency_texture[13][37] = 0;	doodle_right_transparency_texture[13][38] = 0;	doodle_right_transparency_texture[13][39] = 0;	doodle_right_transparency_texture[13][40] = 0;	doodle_right_transparency_texture[13][41] = 0;	doodle_right_transparency_texture[13][42] = 0;	doodle_right_transparency_texture[13][43] = 0;	doodle_right_transparency_texture[13][44] = 0;	doodle_right_transparency_texture[13][45] = 0;	doodle_right_transparency_texture[13][46] = 0;	doodle_right_transparency_texture[13][47] = 0;	doodle_right_transparency_texture[13][48] = 1;	doodle_right_transparency_texture[13][49] = 1;	doodle_right_transparency_texture[13][50] = 1;	doodle_right_transparency_texture[13][51] = 1;	doodle_right_transparency_texture[13][52] = 1;	doodle_right_transparency_texture[13][53] = 1;	doodle_right_transparency_texture[13][54] = 1;	doodle_right_transparency_texture[13][55] = 1;	doodle_right_transparency_texture[13][56] = 1;	doodle_right_transparency_texture[13][57] = 1;	doodle_right_transparency_texture[13][58] = 1;	doodle_right_transparency_texture[13][59] = 1;	doodle_right_transparency_texture[13][60] = 1;	doodle_right_transparency_texture[13][61] = 1;	doodle_right_transparency_texture[13][62] = 1;	doodle_right_transparency_texture[13][63] = 1;	doodle_right_transparency_texture[13][64] = 1;	doodle_right_transparency_texture[13][65] = 1;	doodle_right_transparency_texture[13][66] = 1;	doodle_right_transparency_texture[13][67] = 1;	doodle_right_transparency_texture[13][68] = 1;	doodle_right_transparency_texture[13][69] = 1;	doodle_right_transparency_texture[13][70] = 1;	doodle_right_transparency_texture[13][71] = 1;	doodle_right_transparency_texture[13][72] = 1;	doodle_right_transparency_texture[13][73] = 1;	doodle_right_transparency_texture[13][74] = 1;	doodle_right_transparency_texture[13][75] = 1;	doodle_right_transparency_texture[13][76] = 1;	doodle_right_transparency_texture[13][77] = 1;	doodle_right_transparency_texture[13][78] = 1;	doodle_right_transparency_texture[13][79] = 1;	doodle_right_transparency_texture[14][0] = 1;	doodle_right_transparency_texture[14][1] = 1;	doodle_right_transparency_texture[14][2] = 1;	doodle_right_transparency_texture[14][3] = 1;	doodle_right_transparency_texture[14][4] = 1;	doodle_right_transparency_texture[14][5] = 1;	doodle_right_transparency_texture[14][6] = 1;	doodle_right_transparency_texture[14][7] = 1;	doodle_right_transparency_texture[14][8] = 0;	doodle_right_transparency_texture[14][9] = 0;	doodle_right_transparency_texture[14][10] = 0;	doodle_right_transparency_texture[14][11] = 0;	doodle_right_transparency_texture[14][12] = 0;	doodle_right_transparency_texture[14][13] = 0;	doodle_right_transparency_texture[14][14] = 0;	doodle_right_transparency_texture[14][15] = 0;	doodle_right_transparency_texture[14][16] = 0;	doodle_right_transparency_texture[14][17] = 0;	doodle_right_transparency_texture[14][18] = 0;	doodle_right_transparency_texture[14][19] = 0;	doodle_right_transparency_texture[14][20] = 0;	doodle_right_transparency_texture[14][21] = 0;	doodle_right_transparency_texture[14][22] = 0;	doodle_right_transparency_texture[14][23] = 0;	doodle_right_transparency_texture[14][24] = 0;	doodle_right_transparency_texture[14][25] = 0;	doodle_right_transparency_texture[14][26] = 0;	doodle_right_transparency_texture[14][27] = 0;	doodle_right_transparency_texture[14][28] = 0;	doodle_right_transparency_texture[14][29] = 0;	doodle_right_transparency_texture[14][30] = 0;	doodle_right_transparency_texture[14][31] = 0;	doodle_right_transparency_texture[14][32] = 0;	doodle_right_transparency_texture[14][33] = 0;	doodle_right_transparency_texture[14][34] = 0;	doodle_right_transparency_texture[14][35] = 0;	doodle_right_transparency_texture[14][36] = 0;	doodle_right_transparency_texture[14][37] = 0;	doodle_right_transparency_texture[14][38] = 0;	doodle_right_transparency_texture[14][39] = 0;	doodle_right_transparency_texture[14][40] = 0;	doodle_right_transparency_texture[14][41] = 0;	doodle_right_transparency_texture[14][42] = 0;	doodle_right_transparency_texture[14][43] = 0;	doodle_right_transparency_texture[14][44] = 0;	doodle_right_transparency_texture[14][45] = 0;	doodle_right_transparency_texture[14][46] = 0;	doodle_right_transparency_texture[14][47] = 0;	doodle_right_transparency_texture[14][48] = 1;	doodle_right_transparency_texture[14][49] = 1;	doodle_right_transparency_texture[14][50] = 1;	doodle_right_transparency_texture[14][51] = 1;	doodle_right_transparency_texture[14][52] = 1;	doodle_right_transparency_texture[14][53] = 1;	doodle_right_transparency_texture[14][54] = 1;	doodle_right_transparency_texture[14][55] = 1;	doodle_right_transparency_texture[14][56] = 1;	doodle_right_transparency_texture[14][57] = 1;	doodle_right_transparency_texture[14][58] = 1;	doodle_right_transparency_texture[14][59] = 1;	doodle_right_transparency_texture[14][60] = 1;	doodle_right_transparency_texture[14][61] = 1;	doodle_right_transparency_texture[14][62] = 1;	doodle_right_transparency_texture[14][63] = 1;	doodle_right_transparency_texture[14][64] = 1;	doodle_right_transparency_texture[14][65] = 1;	doodle_right_transparency_texture[14][66] = 1;	doodle_right_transparency_texture[14][67] = 1;	doodle_right_transparency_texture[14][68] = 1;	doodle_right_transparency_texture[14][69] = 1;	doodle_right_transparency_texture[14][70] = 1;	doodle_right_transparency_texture[14][71] = 1;	doodle_right_transparency_texture[14][72] = 1;	doodle_right_transparency_texture[14][73] = 1;	doodle_right_transparency_texture[14][74] = 1;	doodle_right_transparency_texture[14][75] = 1;	doodle_right_transparency_texture[14][76] = 1;	doodle_right_transparency_texture[14][77] = 1;	doodle_right_transparency_texture[14][78] = 1;	doodle_right_transparency_texture[14][79] = 1;	doodle_right_transparency_texture[15][0] = 1;	doodle_right_transparency_texture[15][1] = 1;	doodle_right_transparency_texture[15][2] = 1;	doodle_right_transparency_texture[15][3] = 1;	doodle_right_transparency_texture[15][4] = 1;	doodle_right_transparency_texture[15][5] = 1;	doodle_right_transparency_texture[15][6] = 1;	doodle_right_transparency_texture[15][7] = 1;	doodle_right_transparency_texture[15][8] = 0;	doodle_right_transparency_texture[15][9] = 0;	doodle_right_transparency_texture[15][10] = 0;	doodle_right_transparency_texture[15][11] = 0;	doodle_right_transparency_texture[15][12] = 0;	doodle_right_transparency_texture[15][13] = 0;	doodle_right_transparency_texture[15][14] = 0;	doodle_right_transparency_texture[15][15] = 0;	doodle_right_transparency_texture[15][16] = 0;	doodle_right_transparency_texture[15][17] = 0;	doodle_right_transparency_texture[15][18] = 0;	doodle_right_transparency_texture[15][19] = 0;	doodle_right_transparency_texture[15][20] = 0;	doodle_right_transparency_texture[15][21] = 0;	doodle_right_transparency_texture[15][22] = 0;	doodle_right_transparency_texture[15][23] = 0;	doodle_right_transparency_texture[15][24] = 0;	doodle_right_transparency_texture[15][25] = 0;	doodle_right_transparency_texture[15][26] = 0;	doodle_right_transparency_texture[15][27] = 0;	doodle_right_transparency_texture[15][28] = 0;	doodle_right_transparency_texture[15][29] = 0;	doodle_right_transparency_texture[15][30] = 0;	doodle_right_transparency_texture[15][31] = 0;	doodle_right_transparency_texture[15][32] = 0;	doodle_right_transparency_texture[15][33] = 0;	doodle_right_transparency_texture[15][34] = 0;	doodle_right_transparency_texture[15][35] = 0;	doodle_right_transparency_texture[15][36] = 0;	doodle_right_transparency_texture[15][37] = 0;	doodle_right_transparency_texture[15][38] = 0;	doodle_right_transparency_texture[15][39] = 0;	doodle_right_transparency_texture[15][40] = 0;	doodle_right_transparency_texture[15][41] = 0;	doodle_right_transparency_texture[15][42] = 0;	doodle_right_transparency_texture[15][43] = 0;	doodle_right_transparency_texture[15][44] = 0;	doodle_right_transparency_texture[15][45] = 0;	doodle_right_transparency_texture[15][46] = 0;	doodle_right_transparency_texture[15][47] = 0;	doodle_right_transparency_texture[15][48] = 1;	doodle_right_transparency_texture[15][49] = 1;	doodle_right_transparency_texture[15][50] = 1;	doodle_right_transparency_texture[15][51] = 1;	doodle_right_transparency_texture[15][52] = 1;	doodle_right_transparency_texture[15][53] = 1;	doodle_right_transparency_texture[15][54] = 1;	doodle_right_transparency_texture[15][55] = 1;	doodle_right_transparency_texture[15][56] = 1;	doodle_right_transparency_texture[15][57] = 1;	doodle_right_transparency_texture[15][58] = 1;	doodle_right_transparency_texture[15][59] = 1;	doodle_right_transparency_texture[15][60] = 1;	doodle_right_transparency_texture[15][61] = 1;	doodle_right_transparency_texture[15][62] = 1;	doodle_right_transparency_texture[15][63] = 1;	doodle_right_transparency_texture[15][64] = 1;	doodle_right_transparency_texture[15][65] = 1;	doodle_right_transparency_texture[15][66] = 1;	doodle_right_transparency_texture[15][67] = 1;	doodle_right_transparency_texture[15][68] = 1;	doodle_right_transparency_texture[15][69] = 1;	doodle_right_transparency_texture[15][70] = 1;	doodle_right_transparency_texture[15][71] = 1;	doodle_right_transparency_texture[15][72] = 1;	doodle_right_transparency_texture[15][73] = 1;	doodle_right_transparency_texture[15][74] = 1;	doodle_right_transparency_texture[15][75] = 1;	doodle_right_transparency_texture[15][76] = 1;	doodle_right_transparency_texture[15][77] = 1;	doodle_right_transparency_texture[15][78] = 1;	doodle_right_transparency_texture[15][79] = 1;	doodle_right_transparency_texture[16][0] = 1;	doodle_right_transparency_texture[16][1] = 1;	doodle_right_transparency_texture[16][2] = 1;	doodle_right_transparency_texture[16][3] = 1;	doodle_right_transparency_texture[16][4] = 0;	doodle_right_transparency_texture[16][5] = 0;	doodle_right_transparency_texture[16][6] = 0;	doodle_right_transparency_texture[16][7] = 0;	doodle_right_transparency_texture[16][8] = 0;	doodle_right_transparency_texture[16][9] = 0;	doodle_right_transparency_texture[16][10] = 0;	doodle_right_transparency_texture[16][11] = 0;	doodle_right_transparency_texture[16][12] = 0;	doodle_right_transparency_texture[16][13] = 0;	doodle_right_transparency_texture[16][14] = 0;	doodle_right_transparency_texture[16][15] = 0;	doodle_right_transparency_texture[16][16] = 0;	doodle_right_transparency_texture[16][17] = 0;	doodle_right_transparency_texture[16][18] = 0;	doodle_right_transparency_texture[16][19] = 0;	doodle_right_transparency_texture[16][20] = 0;	doodle_right_transparency_texture[16][21] = 0;	doodle_right_transparency_texture[16][22] = 0;	doodle_right_transparency_texture[16][23] = 0;	doodle_right_transparency_texture[16][24] = 0;	doodle_right_transparency_texture[16][25] = 0;	doodle_right_transparency_texture[16][26] = 0;	doodle_right_transparency_texture[16][27] = 0;	doodle_right_transparency_texture[16][28] = 0;	doodle_right_transparency_texture[16][29] = 0;	doodle_right_transparency_texture[16][30] = 0;	doodle_right_transparency_texture[16][31] = 0;	doodle_right_transparency_texture[16][32] = 0;	doodle_right_transparency_texture[16][33] = 0;	doodle_right_transparency_texture[16][34] = 0;	doodle_right_transparency_texture[16][35] = 0;	doodle_right_transparency_texture[16][36] = 0;	doodle_right_transparency_texture[16][37] = 0;	doodle_right_transparency_texture[16][38] = 0;	doodle_right_transparency_texture[16][39] = 0;	doodle_right_transparency_texture[16][40] = 0;	doodle_right_transparency_texture[16][41] = 0;	doodle_right_transparency_texture[16][42] = 0;	doodle_right_transparency_texture[16][43] = 0;	doodle_right_transparency_texture[16][44] = 0;	doodle_right_transparency_texture[16][45] = 0;	doodle_right_transparency_texture[16][46] = 0;	doodle_right_transparency_texture[16][47] = 0;	doodle_right_transparency_texture[16][48] = 0;	doodle_right_transparency_texture[16][49] = 0;	doodle_right_transparency_texture[16][50] = 0;	doodle_right_transparency_texture[16][51] = 0;	doodle_right_transparency_texture[16][52] = 1;	doodle_right_transparency_texture[16][53] = 1;	doodle_right_transparency_texture[16][54] = 1;	doodle_right_transparency_texture[16][55] = 1;	doodle_right_transparency_texture[16][56] = 1;	doodle_right_transparency_texture[16][57] = 1;	doodle_right_transparency_texture[16][58] = 1;	doodle_right_transparency_texture[16][59] = 1;	doodle_right_transparency_texture[16][60] = 1;	doodle_right_transparency_texture[16][61] = 1;	doodle_right_transparency_texture[16][62] = 1;	doodle_right_transparency_texture[16][63] = 1;	doodle_right_transparency_texture[16][64] = 1;	doodle_right_transparency_texture[16][65] = 1;	doodle_right_transparency_texture[16][66] = 1;	doodle_right_transparency_texture[16][67] = 1;	doodle_right_transparency_texture[16][68] = 1;	doodle_right_transparency_texture[16][69] = 1;	doodle_right_transparency_texture[16][70] = 1;	doodle_right_transparency_texture[16][71] = 1;	doodle_right_transparency_texture[16][72] = 1;	doodle_right_transparency_texture[16][73] = 1;	doodle_right_transparency_texture[16][74] = 1;	doodle_right_transparency_texture[16][75] = 1;	doodle_right_transparency_texture[16][76] = 1;	doodle_right_transparency_texture[16][77] = 1;	doodle_right_transparency_texture[16][78] = 1;	doodle_right_transparency_texture[16][79] = 1;	doodle_right_transparency_texture[17][0] = 1;	doodle_right_transparency_texture[17][1] = 1;	doodle_right_transparency_texture[17][2] = 1;	doodle_right_transparency_texture[17][3] = 1;	doodle_right_transparency_texture[17][4] = 0;	doodle_right_transparency_texture[17][5] = 0;	doodle_right_transparency_texture[17][6] = 0;	doodle_right_transparency_texture[17][7] = 0;	doodle_right_transparency_texture[17][8] = 0;	doodle_right_transparency_texture[17][9] = 0;	doodle_right_transparency_texture[17][10] = 0;	doodle_right_transparency_texture[17][11] = 0;	doodle_right_transparency_texture[17][12] = 0;	doodle_right_transparency_texture[17][13] = 0;	doodle_right_transparency_texture[17][14] = 0;	doodle_right_transparency_texture[17][15] = 0;	doodle_right_transparency_texture[17][16] = 0;	doodle_right_transparency_texture[17][17] = 0;	doodle_right_transparency_texture[17][18] = 0;	doodle_right_transparency_texture[17][19] = 0;	doodle_right_transparency_texture[17][20] = 0;	doodle_right_transparency_texture[17][21] = 0;	doodle_right_transparency_texture[17][22] = 0;	doodle_right_transparency_texture[17][23] = 0;	doodle_right_transparency_texture[17][24] = 0;	doodle_right_transparency_texture[17][25] = 0;	doodle_right_transparency_texture[17][26] = 0;	doodle_right_transparency_texture[17][27] = 0;	doodle_right_transparency_texture[17][28] = 0;	doodle_right_transparency_texture[17][29] = 0;	doodle_right_transparency_texture[17][30] = 0;	doodle_right_transparency_texture[17][31] = 0;	doodle_right_transparency_texture[17][32] = 0;	doodle_right_transparency_texture[17][33] = 0;	doodle_right_transparency_texture[17][34] = 0;	doodle_right_transparency_texture[17][35] = 0;	doodle_right_transparency_texture[17][36] = 0;	doodle_right_transparency_texture[17][37] = 0;	doodle_right_transparency_texture[17][38] = 0;	doodle_right_transparency_texture[17][39] = 0;	doodle_right_transparency_texture[17][40] = 0;	doodle_right_transparency_texture[17][41] = 0;	doodle_right_transparency_texture[17][42] = 0;	doodle_right_transparency_texture[17][43] = 0;	doodle_right_transparency_texture[17][44] = 0;	doodle_right_transparency_texture[17][45] = 0;	doodle_right_transparency_texture[17][46] = 0;	doodle_right_transparency_texture[17][47] = 0;	doodle_right_transparency_texture[17][48] = 0;	doodle_right_transparency_texture[17][49] = 0;	doodle_right_transparency_texture[17][50] = 0;	doodle_right_transparency_texture[17][51] = 0;	doodle_right_transparency_texture[17][52] = 1;	doodle_right_transparency_texture[17][53] = 1;	doodle_right_transparency_texture[17][54] = 1;	doodle_right_transparency_texture[17][55] = 1;	doodle_right_transparency_texture[17][56] = 1;	doodle_right_transparency_texture[17][57] = 1;	doodle_right_transparency_texture[17][58] = 1;	doodle_right_transparency_texture[17][59] = 1;	doodle_right_transparency_texture[17][60] = 1;	doodle_right_transparency_texture[17][61] = 1;	doodle_right_transparency_texture[17][62] = 1;	doodle_right_transparency_texture[17][63] = 1;	doodle_right_transparency_texture[17][64] = 1;	doodle_right_transparency_texture[17][65] = 1;	doodle_right_transparency_texture[17][66] = 1;	doodle_right_transparency_texture[17][67] = 1;	doodle_right_transparency_texture[17][68] = 1;	doodle_right_transparency_texture[17][69] = 1;	doodle_right_transparency_texture[17][70] = 1;	doodle_right_transparency_texture[17][71] = 1;	doodle_right_transparency_texture[17][72] = 1;	doodle_right_transparency_texture[17][73] = 1;	doodle_right_transparency_texture[17][74] = 1;	doodle_right_transparency_texture[17][75] = 1;	doodle_right_transparency_texture[17][76] = 1;	doodle_right_transparency_texture[17][77] = 1;	doodle_right_transparency_texture[17][78] = 1;	doodle_right_transparency_texture[17][79] = 1;	doodle_right_transparency_texture[18][0] = 1;	doodle_right_transparency_texture[18][1] = 1;	doodle_right_transparency_texture[18][2] = 1;	doodle_right_transparency_texture[18][3] = 1;	doodle_right_transparency_texture[18][4] = 0;	doodle_right_transparency_texture[18][5] = 0;	doodle_right_transparency_texture[18][6] = 0;	doodle_right_transparency_texture[18][7] = 0;	doodle_right_transparency_texture[18][8] = 0;	doodle_right_transparency_texture[18][9] = 0;	doodle_right_transparency_texture[18][10] = 0;	doodle_right_transparency_texture[18][11] = 0;	doodle_right_transparency_texture[18][12] = 0;	doodle_right_transparency_texture[18][13] = 0;	doodle_right_transparency_texture[18][14] = 0;	doodle_right_transparency_texture[18][15] = 0;	doodle_right_transparency_texture[18][16] = 0;	doodle_right_transparency_texture[18][17] = 0;	doodle_right_transparency_texture[18][18] = 0;	doodle_right_transparency_texture[18][19] = 0;	doodle_right_transparency_texture[18][20] = 0;	doodle_right_transparency_texture[18][21] = 0;	doodle_right_transparency_texture[18][22] = 0;	doodle_right_transparency_texture[18][23] = 0;	doodle_right_transparency_texture[18][24] = 0;	doodle_right_transparency_texture[18][25] = 0;	doodle_right_transparency_texture[18][26] = 0;	doodle_right_transparency_texture[18][27] = 0;	doodle_right_transparency_texture[18][28] = 0;	doodle_right_transparency_texture[18][29] = 0;	doodle_right_transparency_texture[18][30] = 0;	doodle_right_transparency_texture[18][31] = 0;	doodle_right_transparency_texture[18][32] = 0;	doodle_right_transparency_texture[18][33] = 0;	doodle_right_transparency_texture[18][34] = 0;	doodle_right_transparency_texture[18][35] = 0;	doodle_right_transparency_texture[18][36] = 0;	doodle_right_transparency_texture[18][37] = 0;	doodle_right_transparency_texture[18][38] = 0;	doodle_right_transparency_texture[18][39] = 0;	doodle_right_transparency_texture[18][40] = 0;	doodle_right_transparency_texture[18][41] = 0;	doodle_right_transparency_texture[18][42] = 0;	doodle_right_transparency_texture[18][43] = 0;	doodle_right_transparency_texture[18][44] = 0;	doodle_right_transparency_texture[18][45] = 0;	doodle_right_transparency_texture[18][46] = 0;	doodle_right_transparency_texture[18][47] = 0;	doodle_right_transparency_texture[18][48] = 0;	doodle_right_transparency_texture[18][49] = 0;	doodle_right_transparency_texture[18][50] = 0;	doodle_right_transparency_texture[18][51] = 0;	doodle_right_transparency_texture[18][52] = 1;	doodle_right_transparency_texture[18][53] = 1;	doodle_right_transparency_texture[18][54] = 1;	doodle_right_transparency_texture[18][55] = 1;	doodle_right_transparency_texture[18][56] = 1;	doodle_right_transparency_texture[18][57] = 1;	doodle_right_transparency_texture[18][58] = 1;	doodle_right_transparency_texture[18][59] = 1;	doodle_right_transparency_texture[18][60] = 1;	doodle_right_transparency_texture[18][61] = 1;	doodle_right_transparency_texture[18][62] = 1;	doodle_right_transparency_texture[18][63] = 1;	doodle_right_transparency_texture[18][64] = 1;	doodle_right_transparency_texture[18][65] = 1;	doodle_right_transparency_texture[18][66] = 1;	doodle_right_transparency_texture[18][67] = 1;	doodle_right_transparency_texture[18][68] = 1;	doodle_right_transparency_texture[18][69] = 1;	doodle_right_transparency_texture[18][70] = 1;	doodle_right_transparency_texture[18][71] = 1;	doodle_right_transparency_texture[18][72] = 1;	doodle_right_transparency_texture[18][73] = 1;	doodle_right_transparency_texture[18][74] = 1;	doodle_right_transparency_texture[18][75] = 1;	doodle_right_transparency_texture[18][76] = 1;	doodle_right_transparency_texture[18][77] = 1;	doodle_right_transparency_texture[18][78] = 1;	doodle_right_transparency_texture[18][79] = 1;	doodle_right_transparency_texture[19][0] = 1;	doodle_right_transparency_texture[19][1] = 1;	doodle_right_transparency_texture[19][2] = 1;	doodle_right_transparency_texture[19][3] = 1;	doodle_right_transparency_texture[19][4] = 0;	doodle_right_transparency_texture[19][5] = 0;	doodle_right_transparency_texture[19][6] = 0;	doodle_right_transparency_texture[19][7] = 0;	doodle_right_transparency_texture[19][8] = 0;	doodle_right_transparency_texture[19][9] = 0;	doodle_right_transparency_texture[19][10] = 0;	doodle_right_transparency_texture[19][11] = 0;	doodle_right_transparency_texture[19][12] = 0;	doodle_right_transparency_texture[19][13] = 0;	doodle_right_transparency_texture[19][14] = 0;	doodle_right_transparency_texture[19][15] = 0;	doodle_right_transparency_texture[19][16] = 0;	doodle_right_transparency_texture[19][17] = 0;	doodle_right_transparency_texture[19][18] = 0;	doodle_right_transparency_texture[19][19] = 0;	doodle_right_transparency_texture[19][20] = 0;	doodle_right_transparency_texture[19][21] = 0;	doodle_right_transparency_texture[19][22] = 0;	doodle_right_transparency_texture[19][23] = 0;	doodle_right_transparency_texture[19][24] = 0;	doodle_right_transparency_texture[19][25] = 0;	doodle_right_transparency_texture[19][26] = 0;	doodle_right_transparency_texture[19][27] = 0;	doodle_right_transparency_texture[19][28] = 0;	doodle_right_transparency_texture[19][29] = 0;	doodle_right_transparency_texture[19][30] = 0;	doodle_right_transparency_texture[19][31] = 0;	doodle_right_transparency_texture[19][32] = 0;	doodle_right_transparency_texture[19][33] = 0;	doodle_right_transparency_texture[19][34] = 0;	doodle_right_transparency_texture[19][35] = 0;	doodle_right_transparency_texture[19][36] = 0;	doodle_right_transparency_texture[19][37] = 0;	doodle_right_transparency_texture[19][38] = 0;	doodle_right_transparency_texture[19][39] = 0;	doodle_right_transparency_texture[19][40] = 0;	doodle_right_transparency_texture[19][41] = 0;	doodle_right_transparency_texture[19][42] = 0;	doodle_right_transparency_texture[19][43] = 0;	doodle_right_transparency_texture[19][44] = 0;	doodle_right_transparency_texture[19][45] = 0;	doodle_right_transparency_texture[19][46] = 0;	doodle_right_transparency_texture[19][47] = 0;	doodle_right_transparency_texture[19][48] = 0;	doodle_right_transparency_texture[19][49] = 0;	doodle_right_transparency_texture[19][50] = 0;	doodle_right_transparency_texture[19][51] = 0;	doodle_right_transparency_texture[19][52] = 1;	doodle_right_transparency_texture[19][53] = 1;	doodle_right_transparency_texture[19][54] = 1;	doodle_right_transparency_texture[19][55] = 1;	doodle_right_transparency_texture[19][56] = 1;	doodle_right_transparency_texture[19][57] = 1;	doodle_right_transparency_texture[19][58] = 1;	doodle_right_transparency_texture[19][59] = 1;	doodle_right_transparency_texture[19][60] = 1;	doodle_right_transparency_texture[19][61] = 1;	doodle_right_transparency_texture[19][62] = 1;	doodle_right_transparency_texture[19][63] = 1;	doodle_right_transparency_texture[19][64] = 1;	doodle_right_transparency_texture[19][65] = 1;	doodle_right_transparency_texture[19][66] = 1;	doodle_right_transparency_texture[19][67] = 1;	doodle_right_transparency_texture[19][68] = 1;	doodle_right_transparency_texture[19][69] = 1;	doodle_right_transparency_texture[19][70] = 1;	doodle_right_transparency_texture[19][71] = 1;	doodle_right_transparency_texture[19][72] = 1;	doodle_right_transparency_texture[19][73] = 1;	doodle_right_transparency_texture[19][74] = 1;	doodle_right_transparency_texture[19][75] = 1;	doodle_right_transparency_texture[19][76] = 1;	doodle_right_transparency_texture[19][77] = 1;	doodle_right_transparency_texture[19][78] = 1;	doodle_right_transparency_texture[19][79] = 1;	doodle_right_transparency_texture[20][0] = 1;	doodle_right_transparency_texture[20][1] = 1;	doodle_right_transparency_texture[20][2] = 1;	doodle_right_transparency_texture[20][3] = 1;	doodle_right_transparency_texture[20][4] = 0;	doodle_right_transparency_texture[20][5] = 0;	doodle_right_transparency_texture[20][6] = 0;	doodle_right_transparency_texture[20][7] = 0;	doodle_right_transparency_texture[20][8] = 0;	doodle_right_transparency_texture[20][9] = 0;	doodle_right_transparency_texture[20][10] = 0;	doodle_right_transparency_texture[20][11] = 0;	doodle_right_transparency_texture[20][12] = 0;	doodle_right_transparency_texture[20][13] = 0;	doodle_right_transparency_texture[20][14] = 0;	doodle_right_transparency_texture[20][15] = 0;	doodle_right_transparency_texture[20][16] = 0;	doodle_right_transparency_texture[20][17] = 0;	doodle_right_transparency_texture[20][18] = 0;	doodle_right_transparency_texture[20][19] = 0;	doodle_right_transparency_texture[20][20] = 0;	doodle_right_transparency_texture[20][21] = 0;	doodle_right_transparency_texture[20][22] = 0;	doodle_right_transparency_texture[20][23] = 0;	doodle_right_transparency_texture[20][24] = 0;	doodle_right_transparency_texture[20][25] = 0;	doodle_right_transparency_texture[20][26] = 0;	doodle_right_transparency_texture[20][27] = 0;	doodle_right_transparency_texture[20][28] = 0;	doodle_right_transparency_texture[20][29] = 0;	doodle_right_transparency_texture[20][30] = 0;	doodle_right_transparency_texture[20][31] = 0;	doodle_right_transparency_texture[20][32] = 0;	doodle_right_transparency_texture[20][33] = 0;	doodle_right_transparency_texture[20][34] = 0;	doodle_right_transparency_texture[20][35] = 0;	doodle_right_transparency_texture[20][36] = 0;	doodle_right_transparency_texture[20][37] = 0;	doodle_right_transparency_texture[20][38] = 0;	doodle_right_transparency_texture[20][39] = 0;	doodle_right_transparency_texture[20][40] = 0;	doodle_right_transparency_texture[20][41] = 0;	doodle_right_transparency_texture[20][42] = 0;	doodle_right_transparency_texture[20][43] = 0;	doodle_right_transparency_texture[20][44] = 0;	doodle_right_transparency_texture[20][45] = 0;	doodle_right_transparency_texture[20][46] = 0;	doodle_right_transparency_texture[20][47] = 0;	doodle_right_transparency_texture[20][48] = 0;	doodle_right_transparency_texture[20][49] = 0;	doodle_right_transparency_texture[20][50] = 0;	doodle_right_transparency_texture[20][51] = 0;	doodle_right_transparency_texture[20][52] = 1;	doodle_right_transparency_texture[20][53] = 1;	doodle_right_transparency_texture[20][54] = 1;	doodle_right_transparency_texture[20][55] = 1;	doodle_right_transparency_texture[20][56] = 1;	doodle_right_transparency_texture[20][57] = 1;	doodle_right_transparency_texture[20][58] = 1;	doodle_right_transparency_texture[20][59] = 1;	doodle_right_transparency_texture[20][60] = 1;	doodle_right_transparency_texture[20][61] = 1;	doodle_right_transparency_texture[20][62] = 1;	doodle_right_transparency_texture[20][63] = 1;	doodle_right_transparency_texture[20][64] = 1;	doodle_right_transparency_texture[20][65] = 1;	doodle_right_transparency_texture[20][66] = 1;	doodle_right_transparency_texture[20][67] = 1;	doodle_right_transparency_texture[20][68] = 1;	doodle_right_transparency_texture[20][69] = 1;	doodle_right_transparency_texture[20][70] = 1;	doodle_right_transparency_texture[20][71] = 1;	doodle_right_transparency_texture[20][72] = 1;	doodle_right_transparency_texture[20][73] = 1;	doodle_right_transparency_texture[20][74] = 1;	doodle_right_transparency_texture[20][75] = 1;	doodle_right_transparency_texture[20][76] = 1;	doodle_right_transparency_texture[20][77] = 1;	doodle_right_transparency_texture[20][78] = 1;	doodle_right_transparency_texture[20][79] = 1;	doodle_right_transparency_texture[21][0] = 1;	doodle_right_transparency_texture[21][1] = 1;	doodle_right_transparency_texture[21][2] = 1;	doodle_right_transparency_texture[21][3] = 1;	doodle_right_transparency_texture[21][4] = 0;	doodle_right_transparency_texture[21][5] = 0;	doodle_right_transparency_texture[21][6] = 0;	doodle_right_transparency_texture[21][7] = 0;	doodle_right_transparency_texture[21][8] = 0;	doodle_right_transparency_texture[21][9] = 0;	doodle_right_transparency_texture[21][10] = 0;	doodle_right_transparency_texture[21][11] = 0;	doodle_right_transparency_texture[21][12] = 0;	doodle_right_transparency_texture[21][13] = 0;	doodle_right_transparency_texture[21][14] = 0;	doodle_right_transparency_texture[21][15] = 0;	doodle_right_transparency_texture[21][16] = 0;	doodle_right_transparency_texture[21][17] = 0;	doodle_right_transparency_texture[21][18] = 0;	doodle_right_transparency_texture[21][19] = 0;	doodle_right_transparency_texture[21][20] = 0;	doodle_right_transparency_texture[21][21] = 0;	doodle_right_transparency_texture[21][22] = 0;	doodle_right_transparency_texture[21][23] = 0;	doodle_right_transparency_texture[21][24] = 0;	doodle_right_transparency_texture[21][25] = 0;	doodle_right_transparency_texture[21][26] = 0;	doodle_right_transparency_texture[21][27] = 0;	doodle_right_transparency_texture[21][28] = 0;	doodle_right_transparency_texture[21][29] = 0;	doodle_right_transparency_texture[21][30] = 0;	doodle_right_transparency_texture[21][31] = 0;	doodle_right_transparency_texture[21][32] = 0;	doodle_right_transparency_texture[21][33] = 0;	doodle_right_transparency_texture[21][34] = 0;	doodle_right_transparency_texture[21][35] = 0;	doodle_right_transparency_texture[21][36] = 0;	doodle_right_transparency_texture[21][37] = 0;	doodle_right_transparency_texture[21][38] = 0;	doodle_right_transparency_texture[21][39] = 0;	doodle_right_transparency_texture[21][40] = 0;	doodle_right_transparency_texture[21][41] = 0;	doodle_right_transparency_texture[21][42] = 0;	doodle_right_transparency_texture[21][43] = 0;	doodle_right_transparency_texture[21][44] = 0;	doodle_right_transparency_texture[21][45] = 0;	doodle_right_transparency_texture[21][46] = 0;	doodle_right_transparency_texture[21][47] = 0;	doodle_right_transparency_texture[21][48] = 0;	doodle_right_transparency_texture[21][49] = 0;	doodle_right_transparency_texture[21][50] = 0;	doodle_right_transparency_texture[21][51] = 0;	doodle_right_transparency_texture[21][52] = 1;	doodle_right_transparency_texture[21][53] = 1;	doodle_right_transparency_texture[21][54] = 1;	doodle_right_transparency_texture[21][55] = 1;	doodle_right_transparency_texture[21][56] = 1;	doodle_right_transparency_texture[21][57] = 1;	doodle_right_transparency_texture[21][58] = 1;	doodle_right_transparency_texture[21][59] = 1;	doodle_right_transparency_texture[21][60] = 1;	doodle_right_transparency_texture[21][61] = 1;	doodle_right_transparency_texture[21][62] = 1;	doodle_right_transparency_texture[21][63] = 1;	doodle_right_transparency_texture[21][64] = 1;	doodle_right_transparency_texture[21][65] = 1;	doodle_right_transparency_texture[21][66] = 1;	doodle_right_transparency_texture[21][67] = 1;	doodle_right_transparency_texture[21][68] = 1;	doodle_right_transparency_texture[21][69] = 1;	doodle_right_transparency_texture[21][70] = 1;	doodle_right_transparency_texture[21][71] = 1;	doodle_right_transparency_texture[21][72] = 1;	doodle_right_transparency_texture[21][73] = 1;	doodle_right_transparency_texture[21][74] = 1;	doodle_right_transparency_texture[21][75] = 1;	doodle_right_transparency_texture[21][76] = 1;	doodle_right_transparency_texture[21][77] = 1;	doodle_right_transparency_texture[21][78] = 1;	doodle_right_transparency_texture[21][79] = 1;	doodle_right_transparency_texture[22][0] = 1;	doodle_right_transparency_texture[22][1] = 1;	doodle_right_transparency_texture[22][2] = 1;	doodle_right_transparency_texture[22][3] = 1;	doodle_right_transparency_texture[22][4] = 0;	doodle_right_transparency_texture[22][5] = 0;	doodle_right_transparency_texture[22][6] = 0;	doodle_right_transparency_texture[22][7] = 0;	doodle_right_transparency_texture[22][8] = 0;	doodle_right_transparency_texture[22][9] = 0;	doodle_right_transparency_texture[22][10] = 0;	doodle_right_transparency_texture[22][11] = 0;	doodle_right_transparency_texture[22][12] = 0;	doodle_right_transparency_texture[22][13] = 0;	doodle_right_transparency_texture[22][14] = 0;	doodle_right_transparency_texture[22][15] = 0;	doodle_right_transparency_texture[22][16] = 0;	doodle_right_transparency_texture[22][17] = 0;	doodle_right_transparency_texture[22][18] = 0;	doodle_right_transparency_texture[22][19] = 0;	doodle_right_transparency_texture[22][20] = 0;	doodle_right_transparency_texture[22][21] = 0;	doodle_right_transparency_texture[22][22] = 0;	doodle_right_transparency_texture[22][23] = 0;	doodle_right_transparency_texture[22][24] = 0;	doodle_right_transparency_texture[22][25] = 0;	doodle_right_transparency_texture[22][26] = 0;	doodle_right_transparency_texture[22][27] = 0;	doodle_right_transparency_texture[22][28] = 0;	doodle_right_transparency_texture[22][29] = 0;	doodle_right_transparency_texture[22][30] = 0;	doodle_right_transparency_texture[22][31] = 0;	doodle_right_transparency_texture[22][32] = 0;	doodle_right_transparency_texture[22][33] = 0;	doodle_right_transparency_texture[22][34] = 0;	doodle_right_transparency_texture[22][35] = 0;	doodle_right_transparency_texture[22][36] = 0;	doodle_right_transparency_texture[22][37] = 0;	doodle_right_transparency_texture[22][38] = 0;	doodle_right_transparency_texture[22][39] = 0;	doodle_right_transparency_texture[22][40] = 0;	doodle_right_transparency_texture[22][41] = 0;	doodle_right_transparency_texture[22][42] = 0;	doodle_right_transparency_texture[22][43] = 0;	doodle_right_transparency_texture[22][44] = 0;	doodle_right_transparency_texture[22][45] = 0;	doodle_right_transparency_texture[22][46] = 0;	doodle_right_transparency_texture[22][47] = 0;	doodle_right_transparency_texture[22][48] = 0;	doodle_right_transparency_texture[22][49] = 0;	doodle_right_transparency_texture[22][50] = 0;	doodle_right_transparency_texture[22][51] = 0;	doodle_right_transparency_texture[22][52] = 1;	doodle_right_transparency_texture[22][53] = 1;	doodle_right_transparency_texture[22][54] = 1;	doodle_right_transparency_texture[22][55] = 1;	doodle_right_transparency_texture[22][56] = 1;	doodle_right_transparency_texture[22][57] = 1;	doodle_right_transparency_texture[22][58] = 1;	doodle_right_transparency_texture[22][59] = 1;	doodle_right_transparency_texture[22][60] = 1;	doodle_right_transparency_texture[22][61] = 1;	doodle_right_transparency_texture[22][62] = 1;	doodle_right_transparency_texture[22][63] = 1;	doodle_right_transparency_texture[22][64] = 1;	doodle_right_transparency_texture[22][65] = 1;	doodle_right_transparency_texture[22][66] = 1;	doodle_right_transparency_texture[22][67] = 1;	doodle_right_transparency_texture[22][68] = 1;	doodle_right_transparency_texture[22][69] = 1;	doodle_right_transparency_texture[22][70] = 1;	doodle_right_transparency_texture[22][71] = 1;	doodle_right_transparency_texture[22][72] = 1;	doodle_right_transparency_texture[22][73] = 1;	doodle_right_transparency_texture[22][74] = 1;	doodle_right_transparency_texture[22][75] = 1;	doodle_right_transparency_texture[22][76] = 1;	doodle_right_transparency_texture[22][77] = 1;	doodle_right_transparency_texture[22][78] = 1;	doodle_right_transparency_texture[22][79] = 1;	doodle_right_transparency_texture[23][0] = 1;	doodle_right_transparency_texture[23][1] = 1;	doodle_right_transparency_texture[23][2] = 1;	doodle_right_transparency_texture[23][3] = 1;	doodle_right_transparency_texture[23][4] = 0;	doodle_right_transparency_texture[23][5] = 0;	doodle_right_transparency_texture[23][6] = 0;	doodle_right_transparency_texture[23][7] = 0;	doodle_right_transparency_texture[23][8] = 0;	doodle_right_transparency_texture[23][9] = 0;	doodle_right_transparency_texture[23][10] = 0;	doodle_right_transparency_texture[23][11] = 0;	doodle_right_transparency_texture[23][12] = 0;	doodle_right_transparency_texture[23][13] = 0;	doodle_right_transparency_texture[23][14] = 0;	doodle_right_transparency_texture[23][15] = 0;	doodle_right_transparency_texture[23][16] = 0;	doodle_right_transparency_texture[23][17] = 0;	doodle_right_transparency_texture[23][18] = 0;	doodle_right_transparency_texture[23][19] = 0;	doodle_right_transparency_texture[23][20] = 0;	doodle_right_transparency_texture[23][21] = 0;	doodle_right_transparency_texture[23][22] = 0;	doodle_right_transparency_texture[23][23] = 0;	doodle_right_transparency_texture[23][24] = 0;	doodle_right_transparency_texture[23][25] = 0;	doodle_right_transparency_texture[23][26] = 0;	doodle_right_transparency_texture[23][27] = 0;	doodle_right_transparency_texture[23][28] = 0;	doodle_right_transparency_texture[23][29] = 0;	doodle_right_transparency_texture[23][30] = 0;	doodle_right_transparency_texture[23][31] = 0;	doodle_right_transparency_texture[23][32] = 0;	doodle_right_transparency_texture[23][33] = 0;	doodle_right_transparency_texture[23][34] = 0;	doodle_right_transparency_texture[23][35] = 0;	doodle_right_transparency_texture[23][36] = 0;	doodle_right_transparency_texture[23][37] = 0;	doodle_right_transparency_texture[23][38] = 0;	doodle_right_transparency_texture[23][39] = 0;	doodle_right_transparency_texture[23][40] = 0;	doodle_right_transparency_texture[23][41] = 0;	doodle_right_transparency_texture[23][42] = 0;	doodle_right_transparency_texture[23][43] = 0;	doodle_right_transparency_texture[23][44] = 0;	doodle_right_transparency_texture[23][45] = 0;	doodle_right_transparency_texture[23][46] = 0;	doodle_right_transparency_texture[23][47] = 0;	doodle_right_transparency_texture[23][48] = 0;	doodle_right_transparency_texture[23][49] = 0;	doodle_right_transparency_texture[23][50] = 0;	doodle_right_transparency_texture[23][51] = 0;	doodle_right_transparency_texture[23][52] = 1;	doodle_right_transparency_texture[23][53] = 1;	doodle_right_transparency_texture[23][54] = 1;	doodle_right_transparency_texture[23][55] = 1;	doodle_right_transparency_texture[23][56] = 1;	doodle_right_transparency_texture[23][57] = 1;	doodle_right_transparency_texture[23][58] = 1;	doodle_right_transparency_texture[23][59] = 1;	doodle_right_transparency_texture[23][60] = 1;	doodle_right_transparency_texture[23][61] = 1;	doodle_right_transparency_texture[23][62] = 1;	doodle_right_transparency_texture[23][63] = 1;	doodle_right_transparency_texture[23][64] = 1;	doodle_right_transparency_texture[23][65] = 1;	doodle_right_transparency_texture[23][66] = 1;	doodle_right_transparency_texture[23][67] = 1;	doodle_right_transparency_texture[23][68] = 1;	doodle_right_transparency_texture[23][69] = 1;	doodle_right_transparency_texture[23][70] = 1;	doodle_right_transparency_texture[23][71] = 1;	doodle_right_transparency_texture[23][72] = 1;	doodle_right_transparency_texture[23][73] = 1;	doodle_right_transparency_texture[23][74] = 1;	doodle_right_transparency_texture[23][75] = 1;	doodle_right_transparency_texture[23][76] = 1;	doodle_right_transparency_texture[23][77] = 1;	doodle_right_transparency_texture[23][78] = 1;	doodle_right_transparency_texture[23][79] = 1;	doodle_right_transparency_texture[24][0] = 1;	doodle_right_transparency_texture[24][1] = 1;	doodle_right_transparency_texture[24][2] = 1;	doodle_right_transparency_texture[24][3] = 1;	doodle_right_transparency_texture[24][4] = 0;	doodle_right_transparency_texture[24][5] = 0;	doodle_right_transparency_texture[24][6] = 0;	doodle_right_transparency_texture[24][7] = 0;	doodle_right_transparency_texture[24][8] = 0;	doodle_right_transparency_texture[24][9] = 0;	doodle_right_transparency_texture[24][10] = 0;	doodle_right_transparency_texture[24][11] = 0;	doodle_right_transparency_texture[24][12] = 0;	doodle_right_transparency_texture[24][13] = 0;	doodle_right_transparency_texture[24][14] = 0;	doodle_right_transparency_texture[24][15] = 0;	doodle_right_transparency_texture[24][16] = 0;	doodle_right_transparency_texture[24][17] = 0;	doodle_right_transparency_texture[24][18] = 0;	doodle_right_transparency_texture[24][19] = 0;	doodle_right_transparency_texture[24][20] = 0;	doodle_right_transparency_texture[24][21] = 0;	doodle_right_transparency_texture[24][22] = 0;	doodle_right_transparency_texture[24][23] = 0;	doodle_right_transparency_texture[24][24] = 0;	doodle_right_transparency_texture[24][25] = 0;	doodle_right_transparency_texture[24][26] = 0;	doodle_right_transparency_texture[24][27] = 0;	doodle_right_transparency_texture[24][28] = 0;	doodle_right_transparency_texture[24][29] = 0;	doodle_right_transparency_texture[24][30] = 0;	doodle_right_transparency_texture[24][31] = 0;	doodle_right_transparency_texture[24][32] = 0;	doodle_right_transparency_texture[24][33] = 0;	doodle_right_transparency_texture[24][34] = 0;	doodle_right_transparency_texture[24][35] = 0;	doodle_right_transparency_texture[24][36] = 0;	doodle_right_transparency_texture[24][37] = 0;	doodle_right_transparency_texture[24][38] = 0;	doodle_right_transparency_texture[24][39] = 0;	doodle_right_transparency_texture[24][40] = 0;	doodle_right_transparency_texture[24][41] = 0;	doodle_right_transparency_texture[24][42] = 0;	doodle_right_transparency_texture[24][43] = 0;	doodle_right_transparency_texture[24][44] = 0;	doodle_right_transparency_texture[24][45] = 0;	doodle_right_transparency_texture[24][46] = 0;	doodle_right_transparency_texture[24][47] = 0;	doodle_right_transparency_texture[24][48] = 0;	doodle_right_transparency_texture[24][49] = 0;	doodle_right_transparency_texture[24][50] = 0;	doodle_right_transparency_texture[24][51] = 0;	doodle_right_transparency_texture[24][52] = 0;	doodle_right_transparency_texture[24][53] = 0;	doodle_right_transparency_texture[24][54] = 0;	doodle_right_transparency_texture[24][55] = 0;	doodle_right_transparency_texture[24][56] = 0;	doodle_right_transparency_texture[24][57] = 0;	doodle_right_transparency_texture[24][58] = 0;	doodle_right_transparency_texture[24][59] = 0;	doodle_right_transparency_texture[24][60] = 0;	doodle_right_transparency_texture[24][61] = 0;	doodle_right_transparency_texture[24][62] = 0;	doodle_right_transparency_texture[24][63] = 0;	doodle_right_transparency_texture[24][64] = 0;	doodle_right_transparency_texture[24][65] = 0;	doodle_right_transparency_texture[24][66] = 0;	doodle_right_transparency_texture[24][67] = 0;	doodle_right_transparency_texture[24][68] = 0;	doodle_right_transparency_texture[24][69] = 0;	doodle_right_transparency_texture[24][70] = 0;	doodle_right_transparency_texture[24][71] = 0;	doodle_right_transparency_texture[24][72] = 0;	doodle_right_transparency_texture[24][73] = 0;	doodle_right_transparency_texture[24][74] = 0;	doodle_right_transparency_texture[24][75] = 0;	doodle_right_transparency_texture[24][76] = 1;	doodle_right_transparency_texture[24][77] = 1;	doodle_right_transparency_texture[24][78] = 1;	doodle_right_transparency_texture[24][79] = 1;	doodle_right_transparency_texture[25][0] = 1;	doodle_right_transparency_texture[25][1] = 1;	doodle_right_transparency_texture[25][2] = 1;	doodle_right_transparency_texture[25][3] = 1;	doodle_right_transparency_texture[25][4] = 0;	doodle_right_transparency_texture[25][5] = 0;	doodle_right_transparency_texture[25][6] = 0;	doodle_right_transparency_texture[25][7] = 0;	doodle_right_transparency_texture[25][8] = 0;	doodle_right_transparency_texture[25][9] = 0;	doodle_right_transparency_texture[25][10] = 0;	doodle_right_transparency_texture[25][11] = 0;	doodle_right_transparency_texture[25][12] = 0;	doodle_right_transparency_texture[25][13] = 0;	doodle_right_transparency_texture[25][14] = 0;	doodle_right_transparency_texture[25][15] = 0;	doodle_right_transparency_texture[25][16] = 0;	doodle_right_transparency_texture[25][17] = 0;	doodle_right_transparency_texture[25][18] = 0;	doodle_right_transparency_texture[25][19] = 0;	doodle_right_transparency_texture[25][20] = 0;	doodle_right_transparency_texture[25][21] = 0;	doodle_right_transparency_texture[25][22] = 0;	doodle_right_transparency_texture[25][23] = 0;	doodle_right_transparency_texture[25][24] = 0;	doodle_right_transparency_texture[25][25] = 0;	doodle_right_transparency_texture[25][26] = 0;	doodle_right_transparency_texture[25][27] = 0;	doodle_right_transparency_texture[25][28] = 0;	doodle_right_transparency_texture[25][29] = 0;	doodle_right_transparency_texture[25][30] = 0;	doodle_right_transparency_texture[25][31] = 0;	doodle_right_transparency_texture[25][32] = 0;	doodle_right_transparency_texture[25][33] = 0;	doodle_right_transparency_texture[25][34] = 0;	doodle_right_transparency_texture[25][35] = 0;	doodle_right_transparency_texture[25][36] = 0;	doodle_right_transparency_texture[25][37] = 0;	doodle_right_transparency_texture[25][38] = 0;	doodle_right_transparency_texture[25][39] = 0;	doodle_right_transparency_texture[25][40] = 0;	doodle_right_transparency_texture[25][41] = 0;	doodle_right_transparency_texture[25][42] = 0;	doodle_right_transparency_texture[25][43] = 0;	doodle_right_transparency_texture[25][44] = 0;	doodle_right_transparency_texture[25][45] = 0;	doodle_right_transparency_texture[25][46] = 0;	doodle_right_transparency_texture[25][47] = 0;	doodle_right_transparency_texture[25][48] = 0;	doodle_right_transparency_texture[25][49] = 0;	doodle_right_transparency_texture[25][50] = 0;	doodle_right_transparency_texture[25][51] = 0;	doodle_right_transparency_texture[25][52] = 0;	doodle_right_transparency_texture[25][53] = 0;	doodle_right_transparency_texture[25][54] = 0;	doodle_right_transparency_texture[25][55] = 0;	doodle_right_transparency_texture[25][56] = 0;	doodle_right_transparency_texture[25][57] = 0;	doodle_right_transparency_texture[25][58] = 0;	doodle_right_transparency_texture[25][59] = 0;	doodle_right_transparency_texture[25][60] = 0;	doodle_right_transparency_texture[25][61] = 0;	doodle_right_transparency_texture[25][62] = 0;	doodle_right_transparency_texture[25][63] = 0;	doodle_right_transparency_texture[25][64] = 0;	doodle_right_transparency_texture[25][65] = 0;	doodle_right_transparency_texture[25][66] = 0;	doodle_right_transparency_texture[25][67] = 0;	doodle_right_transparency_texture[25][68] = 0;	doodle_right_transparency_texture[25][69] = 0;	doodle_right_transparency_texture[25][70] = 0;	doodle_right_transparency_texture[25][71] = 0;	doodle_right_transparency_texture[25][72] = 0;	doodle_right_transparency_texture[25][73] = 0;	doodle_right_transparency_texture[25][74] = 0;	doodle_right_transparency_texture[25][75] = 0;	doodle_right_transparency_texture[25][76] = 1;	doodle_right_transparency_texture[25][77] = 1;	doodle_right_transparency_texture[25][78] = 1;	doodle_right_transparency_texture[25][79] = 1;	doodle_right_transparency_texture[26][0] = 1;	doodle_right_transparency_texture[26][1] = 1;	doodle_right_transparency_texture[26][2] = 1;	doodle_right_transparency_texture[26][3] = 1;	doodle_right_transparency_texture[26][4] = 0;	doodle_right_transparency_texture[26][5] = 0;	doodle_right_transparency_texture[26][6] = 0;	doodle_right_transparency_texture[26][7] = 0;	doodle_right_transparency_texture[26][8] = 0;	doodle_right_transparency_texture[26][9] = 0;	doodle_right_transparency_texture[26][10] = 0;	doodle_right_transparency_texture[26][11] = 0;	doodle_right_transparency_texture[26][12] = 0;	doodle_right_transparency_texture[26][13] = 0;	doodle_right_transparency_texture[26][14] = 0;	doodle_right_transparency_texture[26][15] = 0;	doodle_right_transparency_texture[26][16] = 0;	doodle_right_transparency_texture[26][17] = 0;	doodle_right_transparency_texture[26][18] = 0;	doodle_right_transparency_texture[26][19] = 0;	doodle_right_transparency_texture[26][20] = 0;	doodle_right_transparency_texture[26][21] = 0;	doodle_right_transparency_texture[26][22] = 0;	doodle_right_transparency_texture[26][23] = 0;	doodle_right_transparency_texture[26][24] = 0;	doodle_right_transparency_texture[26][25] = 0;	doodle_right_transparency_texture[26][26] = 0;	doodle_right_transparency_texture[26][27] = 0;	doodle_right_transparency_texture[26][28] = 0;	doodle_right_transparency_texture[26][29] = 0;	doodle_right_transparency_texture[26][30] = 0;	doodle_right_transparency_texture[26][31] = 0;	doodle_right_transparency_texture[26][32] = 0;	doodle_right_transparency_texture[26][33] = 0;	doodle_right_transparency_texture[26][34] = 0;	doodle_right_transparency_texture[26][35] = 0;	doodle_right_transparency_texture[26][36] = 0;	doodle_right_transparency_texture[26][37] = 0;	doodle_right_transparency_texture[26][38] = 0;	doodle_right_transparency_texture[26][39] = 0;	doodle_right_transparency_texture[26][40] = 0;	doodle_right_transparency_texture[26][41] = 0;	doodle_right_transparency_texture[26][42] = 0;	doodle_right_transparency_texture[26][43] = 0;	doodle_right_transparency_texture[26][44] = 0;	doodle_right_transparency_texture[26][45] = 0;	doodle_right_transparency_texture[26][46] = 0;	doodle_right_transparency_texture[26][47] = 0;	doodle_right_transparency_texture[26][48] = 0;	doodle_right_transparency_texture[26][49] = 0;	doodle_right_transparency_texture[26][50] = 0;	doodle_right_transparency_texture[26][51] = 0;	doodle_right_transparency_texture[26][52] = 0;	doodle_right_transparency_texture[26][53] = 0;	doodle_right_transparency_texture[26][54] = 0;	doodle_right_transparency_texture[26][55] = 0;	doodle_right_transparency_texture[26][56] = 0;	doodle_right_transparency_texture[26][57] = 0;	doodle_right_transparency_texture[26][58] = 0;	doodle_right_transparency_texture[26][59] = 0;	doodle_right_transparency_texture[26][60] = 0;	doodle_right_transparency_texture[26][61] = 0;	doodle_right_transparency_texture[26][62] = 0;	doodle_right_transparency_texture[26][63] = 0;	doodle_right_transparency_texture[26][64] = 0;	doodle_right_transparency_texture[26][65] = 0;	doodle_right_transparency_texture[26][66] = 0;	doodle_right_transparency_texture[26][67] = 0;	doodle_right_transparency_texture[26][68] = 0;	doodle_right_transparency_texture[26][69] = 0;	doodle_right_transparency_texture[26][70] = 0;	doodle_right_transparency_texture[26][71] = 0;	doodle_right_transparency_texture[26][72] = 0;	doodle_right_transparency_texture[26][73] = 0;	doodle_right_transparency_texture[26][74] = 0;	doodle_right_transparency_texture[26][75] = 0;	doodle_right_transparency_texture[26][76] = 1;	doodle_right_transparency_texture[26][77] = 1;	doodle_right_transparency_texture[26][78] = 1;	doodle_right_transparency_texture[26][79] = 1;	doodle_right_transparency_texture[27][0] = 1;	doodle_right_transparency_texture[27][1] = 1;	doodle_right_transparency_texture[27][2] = 1;	doodle_right_transparency_texture[27][3] = 1;	doodle_right_transparency_texture[27][4] = 0;	doodle_right_transparency_texture[27][5] = 0;	doodle_right_transparency_texture[27][6] = 0;	doodle_right_transparency_texture[27][7] = 0;	doodle_right_transparency_texture[27][8] = 0;	doodle_right_transparency_texture[27][9] = 0;	doodle_right_transparency_texture[27][10] = 0;	doodle_right_transparency_texture[27][11] = 0;	doodle_right_transparency_texture[27][12] = 0;	doodle_right_transparency_texture[27][13] = 0;	doodle_right_transparency_texture[27][14] = 0;	doodle_right_transparency_texture[27][15] = 0;	doodle_right_transparency_texture[27][16] = 0;	doodle_right_transparency_texture[27][17] = 0;	doodle_right_transparency_texture[27][18] = 0;	doodle_right_transparency_texture[27][19] = 0;	doodle_right_transparency_texture[27][20] = 0;	doodle_right_transparency_texture[27][21] = 0;	doodle_right_transparency_texture[27][22] = 0;	doodle_right_transparency_texture[27][23] = 0;	doodle_right_transparency_texture[27][24] = 0;	doodle_right_transparency_texture[27][25] = 0;	doodle_right_transparency_texture[27][26] = 0;	doodle_right_transparency_texture[27][27] = 0;	doodle_right_transparency_texture[27][28] = 0;	doodle_right_transparency_texture[27][29] = 0;	doodle_right_transparency_texture[27][30] = 0;	doodle_right_transparency_texture[27][31] = 0;	doodle_right_transparency_texture[27][32] = 0;	doodle_right_transparency_texture[27][33] = 0;	doodle_right_transparency_texture[27][34] = 0;	doodle_right_transparency_texture[27][35] = 0;	doodle_right_transparency_texture[27][36] = 0;	doodle_right_transparency_texture[27][37] = 0;	doodle_right_transparency_texture[27][38] = 0;	doodle_right_transparency_texture[27][39] = 0;	doodle_right_transparency_texture[27][40] = 0;	doodle_right_transparency_texture[27][41] = 0;	doodle_right_transparency_texture[27][42] = 0;	doodle_right_transparency_texture[27][43] = 0;	doodle_right_transparency_texture[27][44] = 0;	doodle_right_transparency_texture[27][45] = 0;	doodle_right_transparency_texture[27][46] = 0;	doodle_right_transparency_texture[27][47] = 0;	doodle_right_transparency_texture[27][48] = 0;	doodle_right_transparency_texture[27][49] = 0;	doodle_right_transparency_texture[27][50] = 0;	doodle_right_transparency_texture[27][51] = 0;	doodle_right_transparency_texture[27][52] = 0;	doodle_right_transparency_texture[27][53] = 0;	doodle_right_transparency_texture[27][54] = 0;	doodle_right_transparency_texture[27][55] = 0;	doodle_right_transparency_texture[27][56] = 0;	doodle_right_transparency_texture[27][57] = 0;	doodle_right_transparency_texture[27][58] = 0;	doodle_right_transparency_texture[27][59] = 0;	doodle_right_transparency_texture[27][60] = 0;	doodle_right_transparency_texture[27][61] = 0;	doodle_right_transparency_texture[27][62] = 0;	doodle_right_transparency_texture[27][63] = 0;	doodle_right_transparency_texture[27][64] = 0;	doodle_right_transparency_texture[27][65] = 0;	doodle_right_transparency_texture[27][66] = 0;	doodle_right_transparency_texture[27][67] = 0;	doodle_right_transparency_texture[27][68] = 0;	doodle_right_transparency_texture[27][69] = 0;	doodle_right_transparency_texture[27][70] = 0;	doodle_right_transparency_texture[27][71] = 0;	doodle_right_transparency_texture[27][72] = 0;	doodle_right_transparency_texture[27][73] = 0;	doodle_right_transparency_texture[27][74] = 0;	doodle_right_transparency_texture[27][75] = 0;	doodle_right_transparency_texture[27][76] = 1;	doodle_right_transparency_texture[27][77] = 1;	doodle_right_transparency_texture[27][78] = 1;	doodle_right_transparency_texture[27][79] = 1;	doodle_right_transparency_texture[28][0] = 1;	doodle_right_transparency_texture[28][1] = 1;	doodle_right_transparency_texture[28][2] = 1;	doodle_right_transparency_texture[28][3] = 1;	doodle_right_transparency_texture[28][4] = 0;	doodle_right_transparency_texture[28][5] = 0;	doodle_right_transparency_texture[28][6] = 0;	doodle_right_transparency_texture[28][7] = 0;	doodle_right_transparency_texture[28][8] = 0;	doodle_right_transparency_texture[28][9] = 0;	doodle_right_transparency_texture[28][10] = 0;	doodle_right_transparency_texture[28][11] = 0;	doodle_right_transparency_texture[28][12] = 0;	doodle_right_transparency_texture[28][13] = 0;	doodle_right_transparency_texture[28][14] = 0;	doodle_right_transparency_texture[28][15] = 0;	doodle_right_transparency_texture[28][16] = 0;	doodle_right_transparency_texture[28][17] = 0;	doodle_right_transparency_texture[28][18] = 0;	doodle_right_transparency_texture[28][19] = 0;	doodle_right_transparency_texture[28][20] = 0;	doodle_right_transparency_texture[28][21] = 0;	doodle_right_transparency_texture[28][22] = 0;	doodle_right_transparency_texture[28][23] = 0;	doodle_right_transparency_texture[28][24] = 0;	doodle_right_transparency_texture[28][25] = 0;	doodle_right_transparency_texture[28][26] = 0;	doodle_right_transparency_texture[28][27] = 0;	doodle_right_transparency_texture[28][28] = 0;	doodle_right_transparency_texture[28][29] = 0;	doodle_right_transparency_texture[28][30] = 0;	doodle_right_transparency_texture[28][31] = 0;	doodle_right_transparency_texture[28][32] = 0;	doodle_right_transparency_texture[28][33] = 0;	doodle_right_transparency_texture[28][34] = 0;	doodle_right_transparency_texture[28][35] = 0;	doodle_right_transparency_texture[28][36] = 0;	doodle_right_transparency_texture[28][37] = 0;	doodle_right_transparency_texture[28][38] = 0;	doodle_right_transparency_texture[28][39] = 0;	doodle_right_transparency_texture[28][40] = 0;	doodle_right_transparency_texture[28][41] = 0;	doodle_right_transparency_texture[28][42] = 0;	doodle_right_transparency_texture[28][43] = 0;	doodle_right_transparency_texture[28][44] = 0;	doodle_right_transparency_texture[28][45] = 0;	doodle_right_transparency_texture[28][46] = 0;	doodle_right_transparency_texture[28][47] = 0;	doodle_right_transparency_texture[28][48] = 0;	doodle_right_transparency_texture[28][49] = 0;	doodle_right_transparency_texture[28][50] = 0;	doodle_right_transparency_texture[28][51] = 0;	doodle_right_transparency_texture[28][52] = 0;	doodle_right_transparency_texture[28][53] = 0;	doodle_right_transparency_texture[28][54] = 0;	doodle_right_transparency_texture[28][55] = 0;	doodle_right_transparency_texture[28][56] = 0;	doodle_right_transparency_texture[28][57] = 0;	doodle_right_transparency_texture[28][58] = 0;	doodle_right_transparency_texture[28][59] = 0;	doodle_right_transparency_texture[28][60] = 0;	doodle_right_transparency_texture[28][61] = 0;	doodle_right_transparency_texture[28][62] = 0;	doodle_right_transparency_texture[28][63] = 0;	doodle_right_transparency_texture[28][64] = 0;	doodle_right_transparency_texture[28][65] = 0;	doodle_right_transparency_texture[28][66] = 0;	doodle_right_transparency_texture[28][67] = 0;	doodle_right_transparency_texture[28][68] = 0;	doodle_right_transparency_texture[28][69] = 0;	doodle_right_transparency_texture[28][70] = 0;	doodle_right_transparency_texture[28][71] = 0;	doodle_right_transparency_texture[28][72] = 0;	doodle_right_transparency_texture[28][73] = 0;	doodle_right_transparency_texture[28][74] = 0;	doodle_right_transparency_texture[28][75] = 0;	doodle_right_transparency_texture[28][76] = 1;	doodle_right_transparency_texture[28][77] = 1;	doodle_right_transparency_texture[28][78] = 1;	doodle_right_transparency_texture[28][79] = 1;	doodle_right_transparency_texture[29][0] = 1;	doodle_right_transparency_texture[29][1] = 1;	doodle_right_transparency_texture[29][2] = 1;	doodle_right_transparency_texture[29][3] = 1;	doodle_right_transparency_texture[29][4] = 0;	doodle_right_transparency_texture[29][5] = 0;	doodle_right_transparency_texture[29][6] = 0;	doodle_right_transparency_texture[29][7] = 0;	doodle_right_transparency_texture[29][8] = 0;	doodle_right_transparency_texture[29][9] = 0;	doodle_right_transparency_texture[29][10] = 0;	doodle_right_transparency_texture[29][11] = 0;	doodle_right_transparency_texture[29][12] = 0;	doodle_right_transparency_texture[29][13] = 0;	doodle_right_transparency_texture[29][14] = 0;	doodle_right_transparency_texture[29][15] = 0;	doodle_right_transparency_texture[29][16] = 0;	doodle_right_transparency_texture[29][17] = 0;	doodle_right_transparency_texture[29][18] = 0;	doodle_right_transparency_texture[29][19] = 0;	doodle_right_transparency_texture[29][20] = 0;	doodle_right_transparency_texture[29][21] = 0;	doodle_right_transparency_texture[29][22] = 0;	doodle_right_transparency_texture[29][23] = 0;	doodle_right_transparency_texture[29][24] = 0;	doodle_right_transparency_texture[29][25] = 0;	doodle_right_transparency_texture[29][26] = 0;	doodle_right_transparency_texture[29][27] = 0;	doodle_right_transparency_texture[29][28] = 0;	doodle_right_transparency_texture[29][29] = 0;	doodle_right_transparency_texture[29][30] = 0;	doodle_right_transparency_texture[29][31] = 0;	doodle_right_transparency_texture[29][32] = 0;	doodle_right_transparency_texture[29][33] = 0;	doodle_right_transparency_texture[29][34] = 0;	doodle_right_transparency_texture[29][35] = 0;	doodle_right_transparency_texture[29][36] = 0;	doodle_right_transparency_texture[29][37] = 0;	doodle_right_transparency_texture[29][38] = 0;	doodle_right_transparency_texture[29][39] = 0;	doodle_right_transparency_texture[29][40] = 0;	doodle_right_transparency_texture[29][41] = 0;	doodle_right_transparency_texture[29][42] = 0;	doodle_right_transparency_texture[29][43] = 0;	doodle_right_transparency_texture[29][44] = 0;	doodle_right_transparency_texture[29][45] = 0;	doodle_right_transparency_texture[29][46] = 0;	doodle_right_transparency_texture[29][47] = 0;	doodle_right_transparency_texture[29][48] = 0;	doodle_right_transparency_texture[29][49] = 0;	doodle_right_transparency_texture[29][50] = 0;	doodle_right_transparency_texture[29][51] = 0;	doodle_right_transparency_texture[29][52] = 0;	doodle_right_transparency_texture[29][53] = 0;	doodle_right_transparency_texture[29][54] = 0;	doodle_right_transparency_texture[29][55] = 0;	doodle_right_transparency_texture[29][56] = 0;	doodle_right_transparency_texture[29][57] = 0;	doodle_right_transparency_texture[29][58] = 0;	doodle_right_transparency_texture[29][59] = 0;	doodle_right_transparency_texture[29][60] = 0;	doodle_right_transparency_texture[29][61] = 0;	doodle_right_transparency_texture[29][62] = 0;	doodle_right_transparency_texture[29][63] = 0;	doodle_right_transparency_texture[29][64] = 0;	doodle_right_transparency_texture[29][65] = 0;	doodle_right_transparency_texture[29][66] = 0;	doodle_right_transparency_texture[29][67] = 0;	doodle_right_transparency_texture[29][68] = 0;	doodle_right_transparency_texture[29][69] = 0;	doodle_right_transparency_texture[29][70] = 0;	doodle_right_transparency_texture[29][71] = 0;	doodle_right_transparency_texture[29][72] = 0;	doodle_right_transparency_texture[29][73] = 0;	doodle_right_transparency_texture[29][74] = 0;	doodle_right_transparency_texture[29][75] = 0;	doodle_right_transparency_texture[29][76] = 1;	doodle_right_transparency_texture[29][77] = 1;	doodle_right_transparency_texture[29][78] = 1;	doodle_right_transparency_texture[29][79] = 1;	doodle_right_transparency_texture[30][0] = 1;	doodle_right_transparency_texture[30][1] = 1;	doodle_right_transparency_texture[30][2] = 1;	doodle_right_transparency_texture[30][3] = 1;	doodle_right_transparency_texture[30][4] = 0;	doodle_right_transparency_texture[30][5] = 0;	doodle_right_transparency_texture[30][6] = 0;	doodle_right_transparency_texture[30][7] = 0;	doodle_right_transparency_texture[30][8] = 0;	doodle_right_transparency_texture[30][9] = 0;	doodle_right_transparency_texture[30][10] = 0;	doodle_right_transparency_texture[30][11] = 0;	doodle_right_transparency_texture[30][12] = 0;	doodle_right_transparency_texture[30][13] = 0;	doodle_right_transparency_texture[30][14] = 0;	doodle_right_transparency_texture[30][15] = 0;	doodle_right_transparency_texture[30][16] = 0;	doodle_right_transparency_texture[30][17] = 0;	doodle_right_transparency_texture[30][18] = 0;	doodle_right_transparency_texture[30][19] = 0;	doodle_right_transparency_texture[30][20] = 0;	doodle_right_transparency_texture[30][21] = 0;	doodle_right_transparency_texture[30][22] = 0;	doodle_right_transparency_texture[30][23] = 0;	doodle_right_transparency_texture[30][24] = 0;	doodle_right_transparency_texture[30][25] = 0;	doodle_right_transparency_texture[30][26] = 0;	doodle_right_transparency_texture[30][27] = 0;	doodle_right_transparency_texture[30][28] = 0;	doodle_right_transparency_texture[30][29] = 0;	doodle_right_transparency_texture[30][30] = 0;	doodle_right_transparency_texture[30][31] = 0;	doodle_right_transparency_texture[30][32] = 0;	doodle_right_transparency_texture[30][33] = 0;	doodle_right_transparency_texture[30][34] = 0;	doodle_right_transparency_texture[30][35] = 0;	doodle_right_transparency_texture[30][36] = 0;	doodle_right_transparency_texture[30][37] = 0;	doodle_right_transparency_texture[30][38] = 0;	doodle_right_transparency_texture[30][39] = 0;	doodle_right_transparency_texture[30][40] = 0;	doodle_right_transparency_texture[30][41] = 0;	doodle_right_transparency_texture[30][42] = 0;	doodle_right_transparency_texture[30][43] = 0;	doodle_right_transparency_texture[30][44] = 0;	doodle_right_transparency_texture[30][45] = 0;	doodle_right_transparency_texture[30][46] = 0;	doodle_right_transparency_texture[30][47] = 0;	doodle_right_transparency_texture[30][48] = 0;	doodle_right_transparency_texture[30][49] = 0;	doodle_right_transparency_texture[30][50] = 0;	doodle_right_transparency_texture[30][51] = 0;	doodle_right_transparency_texture[30][52] = 0;	doodle_right_transparency_texture[30][53] = 0;	doodle_right_transparency_texture[30][54] = 0;	doodle_right_transparency_texture[30][55] = 0;	doodle_right_transparency_texture[30][56] = 0;	doodle_right_transparency_texture[30][57] = 0;	doodle_right_transparency_texture[30][58] = 0;	doodle_right_transparency_texture[30][59] = 0;	doodle_right_transparency_texture[30][60] = 0;	doodle_right_transparency_texture[30][61] = 0;	doodle_right_transparency_texture[30][62] = 0;	doodle_right_transparency_texture[30][63] = 0;	doodle_right_transparency_texture[30][64] = 0;	doodle_right_transparency_texture[30][65] = 0;	doodle_right_transparency_texture[30][66] = 0;	doodle_right_transparency_texture[30][67] = 0;	doodle_right_transparency_texture[30][68] = 0;	doodle_right_transparency_texture[30][69] = 0;	doodle_right_transparency_texture[30][70] = 0;	doodle_right_transparency_texture[30][71] = 0;	doodle_right_transparency_texture[30][72] = 0;	doodle_right_transparency_texture[30][73] = 0;	doodle_right_transparency_texture[30][74] = 0;	doodle_right_transparency_texture[30][75] = 0;	doodle_right_transparency_texture[30][76] = 1;	doodle_right_transparency_texture[30][77] = 1;	doodle_right_transparency_texture[30][78] = 1;	doodle_right_transparency_texture[30][79] = 1;	doodle_right_transparency_texture[31][0] = 1;	doodle_right_transparency_texture[31][1] = 1;	doodle_right_transparency_texture[31][2] = 1;	doodle_right_transparency_texture[31][3] = 1;	doodle_right_transparency_texture[31][4] = 0;	doodle_right_transparency_texture[31][5] = 0;	doodle_right_transparency_texture[31][6] = 0;	doodle_right_transparency_texture[31][7] = 0;	doodle_right_transparency_texture[31][8] = 0;	doodle_right_transparency_texture[31][9] = 0;	doodle_right_transparency_texture[31][10] = 0;	doodle_right_transparency_texture[31][11] = 0;	doodle_right_transparency_texture[31][12] = 0;	doodle_right_transparency_texture[31][13] = 0;	doodle_right_transparency_texture[31][14] = 0;	doodle_right_transparency_texture[31][15] = 0;	doodle_right_transparency_texture[31][16] = 0;	doodle_right_transparency_texture[31][17] = 0;	doodle_right_transparency_texture[31][18] = 0;	doodle_right_transparency_texture[31][19] = 0;	doodle_right_transparency_texture[31][20] = 0;	doodle_right_transparency_texture[31][21] = 0;	doodle_right_transparency_texture[31][22] = 0;	doodle_right_transparency_texture[31][23] = 0;	doodle_right_transparency_texture[31][24] = 0;	doodle_right_transparency_texture[31][25] = 0;	doodle_right_transparency_texture[31][26] = 0;	doodle_right_transparency_texture[31][27] = 0;	doodle_right_transparency_texture[31][28] = 0;	doodle_right_transparency_texture[31][29] = 0;	doodle_right_transparency_texture[31][30] = 0;	doodle_right_transparency_texture[31][31] = 0;	doodle_right_transparency_texture[31][32] = 0;	doodle_right_transparency_texture[31][33] = 0;	doodle_right_transparency_texture[31][34] = 0;	doodle_right_transparency_texture[31][35] = 0;	doodle_right_transparency_texture[31][36] = 0;	doodle_right_transparency_texture[31][37] = 0;	doodle_right_transparency_texture[31][38] = 0;	doodle_right_transparency_texture[31][39] = 0;	doodle_right_transparency_texture[31][40] = 0;	doodle_right_transparency_texture[31][41] = 0;	doodle_right_transparency_texture[31][42] = 0;	doodle_right_transparency_texture[31][43] = 0;	doodle_right_transparency_texture[31][44] = 0;	doodle_right_transparency_texture[31][45] = 0;	doodle_right_transparency_texture[31][46] = 0;	doodle_right_transparency_texture[31][47] = 0;	doodle_right_transparency_texture[31][48] = 0;	doodle_right_transparency_texture[31][49] = 0;	doodle_right_transparency_texture[31][50] = 0;	doodle_right_transparency_texture[31][51] = 0;	doodle_right_transparency_texture[31][52] = 0;	doodle_right_transparency_texture[31][53] = 0;	doodle_right_transparency_texture[31][54] = 0;	doodle_right_transparency_texture[31][55] = 0;	doodle_right_transparency_texture[31][56] = 0;	doodle_right_transparency_texture[31][57] = 0;	doodle_right_transparency_texture[31][58] = 0;	doodle_right_transparency_texture[31][59] = 0;	doodle_right_transparency_texture[31][60] = 0;	doodle_right_transparency_texture[31][61] = 0;	doodle_right_transparency_texture[31][62] = 0;	doodle_right_transparency_texture[31][63] = 0;	doodle_right_transparency_texture[31][64] = 0;	doodle_right_transparency_texture[31][65] = 0;	doodle_right_transparency_texture[31][66] = 0;	doodle_right_transparency_texture[31][67] = 0;	doodle_right_transparency_texture[31][68] = 0;	doodle_right_transparency_texture[31][69] = 0;	doodle_right_transparency_texture[31][70] = 0;	doodle_right_transparency_texture[31][71] = 0;	doodle_right_transparency_texture[31][72] = 0;	doodle_right_transparency_texture[31][73] = 0;	doodle_right_transparency_texture[31][74] = 0;	doodle_right_transparency_texture[31][75] = 0;	doodle_right_transparency_texture[31][76] = 1;	doodle_right_transparency_texture[31][77] = 1;	doodle_right_transparency_texture[31][78] = 1;	doodle_right_transparency_texture[31][79] = 1;	doodle_right_transparency_texture[32][0] = 1;	doodle_right_transparency_texture[32][1] = 1;	doodle_right_transparency_texture[32][2] = 1;	doodle_right_transparency_texture[32][3] = 1;	doodle_right_transparency_texture[32][4] = 0;	doodle_right_transparency_texture[32][5] = 0;	doodle_right_transparency_texture[32][6] = 0;	doodle_right_transparency_texture[32][7] = 0;	doodle_right_transparency_texture[32][8] = 0;	doodle_right_transparency_texture[32][9] = 0;	doodle_right_transparency_texture[32][10] = 0;	doodle_right_transparency_texture[32][11] = 0;	doodle_right_transparency_texture[32][12] = 0;	doodle_right_transparency_texture[32][13] = 0;	doodle_right_transparency_texture[32][14] = 0;	doodle_right_transparency_texture[32][15] = 0;	doodle_right_transparency_texture[32][16] = 0;	doodle_right_transparency_texture[32][17] = 0;	doodle_right_transparency_texture[32][18] = 0;	doodle_right_transparency_texture[32][19] = 0;	doodle_right_transparency_texture[32][20] = 0;	doodle_right_transparency_texture[32][21] = 0;	doodle_right_transparency_texture[32][22] = 0;	doodle_right_transparency_texture[32][23] = 0;	doodle_right_transparency_texture[32][24] = 0;	doodle_right_transparency_texture[32][25] = 0;	doodle_right_transparency_texture[32][26] = 0;	doodle_right_transparency_texture[32][27] = 0;	doodle_right_transparency_texture[32][28] = 0;	doodle_right_transparency_texture[32][29] = 0;	doodle_right_transparency_texture[32][30] = 0;	doodle_right_transparency_texture[32][31] = 0;	doodle_right_transparency_texture[32][32] = 0;	doodle_right_transparency_texture[32][33] = 0;	doodle_right_transparency_texture[32][34] = 0;	doodle_right_transparency_texture[32][35] = 0;	doodle_right_transparency_texture[32][36] = 0;	doodle_right_transparency_texture[32][37] = 0;	doodle_right_transparency_texture[32][38] = 0;	doodle_right_transparency_texture[32][39] = 0;	doodle_right_transparency_texture[32][40] = 0;	doodle_right_transparency_texture[32][41] = 0;	doodle_right_transparency_texture[32][42] = 0;	doodle_right_transparency_texture[32][43] = 0;	doodle_right_transparency_texture[32][44] = 0;	doodle_right_transparency_texture[32][45] = 0;	doodle_right_transparency_texture[32][46] = 0;	doodle_right_transparency_texture[32][47] = 0;	doodle_right_transparency_texture[32][48] = 0;	doodle_right_transparency_texture[32][49] = 0;	doodle_right_transparency_texture[32][50] = 0;	doodle_right_transparency_texture[32][51] = 0;	doodle_right_transparency_texture[32][52] = 0;	doodle_right_transparency_texture[32][53] = 0;	doodle_right_transparency_texture[32][54] = 0;	doodle_right_transparency_texture[32][55] = 0;	doodle_right_transparency_texture[32][56] = 0;	doodle_right_transparency_texture[32][57] = 0;	doodle_right_transparency_texture[32][58] = 0;	doodle_right_transparency_texture[32][59] = 0;	doodle_right_transparency_texture[32][60] = 0;	doodle_right_transparency_texture[32][61] = 0;	doodle_right_transparency_texture[32][62] = 0;	doodle_right_transparency_texture[32][63] = 0;	doodle_right_transparency_texture[32][64] = 0;	doodle_right_transparency_texture[32][65] = 0;	doodle_right_transparency_texture[32][66] = 0;	doodle_right_transparency_texture[32][67] = 0;	doodle_right_transparency_texture[32][68] = 0;	doodle_right_transparency_texture[32][69] = 0;	doodle_right_transparency_texture[32][70] = 0;	doodle_right_transparency_texture[32][71] = 0;	doodle_right_transparency_texture[32][72] = 0;	doodle_right_transparency_texture[32][73] = 0;	doodle_right_transparency_texture[32][74] = 0;	doodle_right_transparency_texture[32][75] = 0;	doodle_right_transparency_texture[32][76] = 1;	doodle_right_transparency_texture[32][77] = 1;	doodle_right_transparency_texture[32][78] = 1;	doodle_right_transparency_texture[32][79] = 1;	doodle_right_transparency_texture[33][0] = 1;	doodle_right_transparency_texture[33][1] = 1;	doodle_right_transparency_texture[33][2] = 1;	doodle_right_transparency_texture[33][3] = 1;	doodle_right_transparency_texture[33][4] = 0;	doodle_right_transparency_texture[33][5] = 0;	doodle_right_transparency_texture[33][6] = 0;	doodle_right_transparency_texture[33][7] = 0;	doodle_right_transparency_texture[33][8] = 0;	doodle_right_transparency_texture[33][9] = 0;	doodle_right_transparency_texture[33][10] = 0;	doodle_right_transparency_texture[33][11] = 0;	doodle_right_transparency_texture[33][12] = 0;	doodle_right_transparency_texture[33][13] = 0;	doodle_right_transparency_texture[33][14] = 0;	doodle_right_transparency_texture[33][15] = 0;	doodle_right_transparency_texture[33][16] = 0;	doodle_right_transparency_texture[33][17] = 0;	doodle_right_transparency_texture[33][18] = 0;	doodle_right_transparency_texture[33][19] = 0;	doodle_right_transparency_texture[33][20] = 0;	doodle_right_transparency_texture[33][21] = 0;	doodle_right_transparency_texture[33][22] = 0;	doodle_right_transparency_texture[33][23] = 0;	doodle_right_transparency_texture[33][24] = 0;	doodle_right_transparency_texture[33][25] = 0;	doodle_right_transparency_texture[33][26] = 0;	doodle_right_transparency_texture[33][27] = 0;	doodle_right_transparency_texture[33][28] = 0;	doodle_right_transparency_texture[33][29] = 0;	doodle_right_transparency_texture[33][30] = 0;	doodle_right_transparency_texture[33][31] = 0;	doodle_right_transparency_texture[33][32] = 0;	doodle_right_transparency_texture[33][33] = 0;	doodle_right_transparency_texture[33][34] = 0;	doodle_right_transparency_texture[33][35] = 0;	doodle_right_transparency_texture[33][36] = 0;	doodle_right_transparency_texture[33][37] = 0;	doodle_right_transparency_texture[33][38] = 0;	doodle_right_transparency_texture[33][39] = 0;	doodle_right_transparency_texture[33][40] = 0;	doodle_right_transparency_texture[33][41] = 0;	doodle_right_transparency_texture[33][42] = 0;	doodle_right_transparency_texture[33][43] = 0;	doodle_right_transparency_texture[33][44] = 0;	doodle_right_transparency_texture[33][45] = 0;	doodle_right_transparency_texture[33][46] = 0;	doodle_right_transparency_texture[33][47] = 0;	doodle_right_transparency_texture[33][48] = 0;	doodle_right_transparency_texture[33][49] = 0;	doodle_right_transparency_texture[33][50] = 0;	doodle_right_transparency_texture[33][51] = 0;	doodle_right_transparency_texture[33][52] = 0;	doodle_right_transparency_texture[33][53] = 0;	doodle_right_transparency_texture[33][54] = 0;	doodle_right_transparency_texture[33][55] = 0;	doodle_right_transparency_texture[33][56] = 0;	doodle_right_transparency_texture[33][57] = 0;	doodle_right_transparency_texture[33][58] = 0;	doodle_right_transparency_texture[33][59] = 0;	doodle_right_transparency_texture[33][60] = 0;	doodle_right_transparency_texture[33][61] = 0;	doodle_right_transparency_texture[33][62] = 0;	doodle_right_transparency_texture[33][63] = 0;	doodle_right_transparency_texture[33][64] = 0;	doodle_right_transparency_texture[33][65] = 0;	doodle_right_transparency_texture[33][66] = 0;	doodle_right_transparency_texture[33][67] = 0;	doodle_right_transparency_texture[33][68] = 0;	doodle_right_transparency_texture[33][69] = 0;	doodle_right_transparency_texture[33][70] = 0;	doodle_right_transparency_texture[33][71] = 0;	doodle_right_transparency_texture[33][72] = 0;	doodle_right_transparency_texture[33][73] = 0;	doodle_right_transparency_texture[33][74] = 0;	doodle_right_transparency_texture[33][75] = 0;	doodle_right_transparency_texture[33][76] = 1;	doodle_right_transparency_texture[33][77] = 1;	doodle_right_transparency_texture[33][78] = 1;	doodle_right_transparency_texture[33][79] = 1;	doodle_right_transparency_texture[34][0] = 1;	doodle_right_transparency_texture[34][1] = 1;	doodle_right_transparency_texture[34][2] = 1;	doodle_right_transparency_texture[34][3] = 1;	doodle_right_transparency_texture[34][4] = 0;	doodle_right_transparency_texture[34][5] = 0;	doodle_right_transparency_texture[34][6] = 0;	doodle_right_transparency_texture[34][7] = 0;	doodle_right_transparency_texture[34][8] = 0;	doodle_right_transparency_texture[34][9] = 0;	doodle_right_transparency_texture[34][10] = 0;	doodle_right_transparency_texture[34][11] = 0;	doodle_right_transparency_texture[34][12] = 0;	doodle_right_transparency_texture[34][13] = 0;	doodle_right_transparency_texture[34][14] = 0;	doodle_right_transparency_texture[34][15] = 0;	doodle_right_transparency_texture[34][16] = 0;	doodle_right_transparency_texture[34][17] = 0;	doodle_right_transparency_texture[34][18] = 0;	doodle_right_transparency_texture[34][19] = 0;	doodle_right_transparency_texture[34][20] = 0;	doodle_right_transparency_texture[34][21] = 0;	doodle_right_transparency_texture[34][22] = 0;	doodle_right_transparency_texture[34][23] = 0;	doodle_right_transparency_texture[34][24] = 0;	doodle_right_transparency_texture[34][25] = 0;	doodle_right_transparency_texture[34][26] = 0;	doodle_right_transparency_texture[34][27] = 0;	doodle_right_transparency_texture[34][28] = 0;	doodle_right_transparency_texture[34][29] = 0;	doodle_right_transparency_texture[34][30] = 0;	doodle_right_transparency_texture[34][31] = 0;	doodle_right_transparency_texture[34][32] = 0;	doodle_right_transparency_texture[34][33] = 0;	doodle_right_transparency_texture[34][34] = 0;	doodle_right_transparency_texture[34][35] = 0;	doodle_right_transparency_texture[34][36] = 0;	doodle_right_transparency_texture[34][37] = 0;	doodle_right_transparency_texture[34][38] = 0;	doodle_right_transparency_texture[34][39] = 0;	doodle_right_transparency_texture[34][40] = 0;	doodle_right_transparency_texture[34][41] = 0;	doodle_right_transparency_texture[34][42] = 0;	doodle_right_transparency_texture[34][43] = 0;	doodle_right_transparency_texture[34][44] = 0;	doodle_right_transparency_texture[34][45] = 0;	doodle_right_transparency_texture[34][46] = 0;	doodle_right_transparency_texture[34][47] = 0;	doodle_right_transparency_texture[34][48] = 0;	doodle_right_transparency_texture[34][49] = 0;	doodle_right_transparency_texture[34][50] = 0;	doodle_right_transparency_texture[34][51] = 0;	doodle_right_transparency_texture[34][52] = 0;	doodle_right_transparency_texture[34][53] = 0;	doodle_right_transparency_texture[34][54] = 0;	doodle_right_transparency_texture[34][55] = 0;	doodle_right_transparency_texture[34][56] = 0;	doodle_right_transparency_texture[34][57] = 0;	doodle_right_transparency_texture[34][58] = 0;	doodle_right_transparency_texture[34][59] = 0;	doodle_right_transparency_texture[34][60] = 0;	doodle_right_transparency_texture[34][61] = 0;	doodle_right_transparency_texture[34][62] = 0;	doodle_right_transparency_texture[34][63] = 0;	doodle_right_transparency_texture[34][64] = 0;	doodle_right_transparency_texture[34][65] = 0;	doodle_right_transparency_texture[34][66] = 0;	doodle_right_transparency_texture[34][67] = 0;	doodle_right_transparency_texture[34][68] = 0;	doodle_right_transparency_texture[34][69] = 0;	doodle_right_transparency_texture[34][70] = 0;	doodle_right_transparency_texture[34][71] = 0;	doodle_right_transparency_texture[34][72] = 0;	doodle_right_transparency_texture[34][73] = 0;	doodle_right_transparency_texture[34][74] = 0;	doodle_right_transparency_texture[34][75] = 0;	doodle_right_transparency_texture[34][76] = 1;	doodle_right_transparency_texture[34][77] = 1;	doodle_right_transparency_texture[34][78] = 1;	doodle_right_transparency_texture[34][79] = 1;	doodle_right_transparency_texture[35][0] = 1;	doodle_right_transparency_texture[35][1] = 1;	doodle_right_transparency_texture[35][2] = 1;	doodle_right_transparency_texture[35][3] = 1;	doodle_right_transparency_texture[35][4] = 0;	doodle_right_transparency_texture[35][5] = 0;	doodle_right_transparency_texture[35][6] = 0;	doodle_right_transparency_texture[35][7] = 0;	doodle_right_transparency_texture[35][8] = 0;	doodle_right_transparency_texture[35][9] = 0;	doodle_right_transparency_texture[35][10] = 0;	doodle_right_transparency_texture[35][11] = 0;	doodle_right_transparency_texture[35][12] = 0;	doodle_right_transparency_texture[35][13] = 0;	doodle_right_transparency_texture[35][14] = 0;	doodle_right_transparency_texture[35][15] = 0;	doodle_right_transparency_texture[35][16] = 0;	doodle_right_transparency_texture[35][17] = 0;	doodle_right_transparency_texture[35][18] = 0;	doodle_right_transparency_texture[35][19] = 0;	doodle_right_transparency_texture[35][20] = 0;	doodle_right_transparency_texture[35][21] = 0;	doodle_right_transparency_texture[35][22] = 0;	doodle_right_transparency_texture[35][23] = 0;	doodle_right_transparency_texture[35][24] = 0;	doodle_right_transparency_texture[35][25] = 0;	doodle_right_transparency_texture[35][26] = 0;	doodle_right_transparency_texture[35][27] = 0;	doodle_right_transparency_texture[35][28] = 0;	doodle_right_transparency_texture[35][29] = 0;	doodle_right_transparency_texture[35][30] = 0;	doodle_right_transparency_texture[35][31] = 0;	doodle_right_transparency_texture[35][32] = 0;	doodle_right_transparency_texture[35][33] = 0;	doodle_right_transparency_texture[35][34] = 0;	doodle_right_transparency_texture[35][35] = 0;	doodle_right_transparency_texture[35][36] = 0;	doodle_right_transparency_texture[35][37] = 0;	doodle_right_transparency_texture[35][38] = 0;	doodle_right_transparency_texture[35][39] = 0;	doodle_right_transparency_texture[35][40] = 0;	doodle_right_transparency_texture[35][41] = 0;	doodle_right_transparency_texture[35][42] = 0;	doodle_right_transparency_texture[35][43] = 0;	doodle_right_transparency_texture[35][44] = 0;	doodle_right_transparency_texture[35][45] = 0;	doodle_right_transparency_texture[35][46] = 0;	doodle_right_transparency_texture[35][47] = 0;	doodle_right_transparency_texture[35][48] = 0;	doodle_right_transparency_texture[35][49] = 0;	doodle_right_transparency_texture[35][50] = 0;	doodle_right_transparency_texture[35][51] = 0;	doodle_right_transparency_texture[35][52] = 0;	doodle_right_transparency_texture[35][53] = 0;	doodle_right_transparency_texture[35][54] = 0;	doodle_right_transparency_texture[35][55] = 0;	doodle_right_transparency_texture[35][56] = 0;	doodle_right_transparency_texture[35][57] = 0;	doodle_right_transparency_texture[35][58] = 0;	doodle_right_transparency_texture[35][59] = 0;	doodle_right_transparency_texture[35][60] = 0;	doodle_right_transparency_texture[35][61] = 0;	doodle_right_transparency_texture[35][62] = 0;	doodle_right_transparency_texture[35][63] = 0;	doodle_right_transparency_texture[35][64] = 0;	doodle_right_transparency_texture[35][65] = 0;	doodle_right_transparency_texture[35][66] = 0;	doodle_right_transparency_texture[35][67] = 0;	doodle_right_transparency_texture[35][68] = 0;	doodle_right_transparency_texture[35][69] = 0;	doodle_right_transparency_texture[35][70] = 0;	doodle_right_transparency_texture[35][71] = 0;	doodle_right_transparency_texture[35][72] = 0;	doodle_right_transparency_texture[35][73] = 0;	doodle_right_transparency_texture[35][74] = 0;	doodle_right_transparency_texture[35][75] = 0;	doodle_right_transparency_texture[35][76] = 1;	doodle_right_transparency_texture[35][77] = 1;	doodle_right_transparency_texture[35][78] = 1;	doodle_right_transparency_texture[35][79] = 1;	doodle_right_transparency_texture[36][0] = 1;	doodle_right_transparency_texture[36][1] = 1;	doodle_right_transparency_texture[36][2] = 1;	doodle_right_transparency_texture[36][3] = 1;	doodle_right_transparency_texture[36][4] = 0;	doodle_right_transparency_texture[36][5] = 0;	doodle_right_transparency_texture[36][6] = 0;	doodle_right_transparency_texture[36][7] = 0;	doodle_right_transparency_texture[36][8] = 0;	doodle_right_transparency_texture[36][9] = 0;	doodle_right_transparency_texture[36][10] = 0;	doodle_right_transparency_texture[36][11] = 0;	doodle_right_transparency_texture[36][12] = 0;	doodle_right_transparency_texture[36][13] = 0;	doodle_right_transparency_texture[36][14] = 0;	doodle_right_transparency_texture[36][15] = 0;	doodle_right_transparency_texture[36][16] = 0;	doodle_right_transparency_texture[36][17] = 0;	doodle_right_transparency_texture[36][18] = 0;	doodle_right_transparency_texture[36][19] = 0;	doodle_right_transparency_texture[36][20] = 0;	doodle_right_transparency_texture[36][21] = 0;	doodle_right_transparency_texture[36][22] = 0;	doodle_right_transparency_texture[36][23] = 0;	doodle_right_transparency_texture[36][24] = 0;	doodle_right_transparency_texture[36][25] = 0;	doodle_right_transparency_texture[36][26] = 0;	doodle_right_transparency_texture[36][27] = 0;	doodle_right_transparency_texture[36][28] = 0;	doodle_right_transparency_texture[36][29] = 0;	doodle_right_transparency_texture[36][30] = 0;	doodle_right_transparency_texture[36][31] = 0;	doodle_right_transparency_texture[36][32] = 0;	doodle_right_transparency_texture[36][33] = 0;	doodle_right_transparency_texture[36][34] = 0;	doodle_right_transparency_texture[36][35] = 0;	doodle_right_transparency_texture[36][36] = 0;	doodle_right_transparency_texture[36][37] = 0;	doodle_right_transparency_texture[36][38] = 0;	doodle_right_transparency_texture[36][39] = 0;	doodle_right_transparency_texture[36][40] = 0;	doodle_right_transparency_texture[36][41] = 0;	doodle_right_transparency_texture[36][42] = 0;	doodle_right_transparency_texture[36][43] = 0;	doodle_right_transparency_texture[36][44] = 0;	doodle_right_transparency_texture[36][45] = 0;	doodle_right_transparency_texture[36][46] = 0;	doodle_right_transparency_texture[36][47] = 0;	doodle_right_transparency_texture[36][48] = 0;	doodle_right_transparency_texture[36][49] = 0;	doodle_right_transparency_texture[36][50] = 0;	doodle_right_transparency_texture[36][51] = 0;	doodle_right_transparency_texture[36][52] = 1;	doodle_right_transparency_texture[36][53] = 1;	doodle_right_transparency_texture[36][54] = 1;	doodle_right_transparency_texture[36][55] = 1;	doodle_right_transparency_texture[36][56] = 1;	doodle_right_transparency_texture[36][57] = 1;	doodle_right_transparency_texture[36][58] = 1;	doodle_right_transparency_texture[36][59] = 1;	doodle_right_transparency_texture[36][60] = 1;	doodle_right_transparency_texture[36][61] = 1;	doodle_right_transparency_texture[36][62] = 1;	doodle_right_transparency_texture[36][63] = 1;	doodle_right_transparency_texture[36][64] = 1;	doodle_right_transparency_texture[36][65] = 1;	doodle_right_transparency_texture[36][66] = 1;	doodle_right_transparency_texture[36][67] = 1;	doodle_right_transparency_texture[36][68] = 1;	doodle_right_transparency_texture[36][69] = 1;	doodle_right_transparency_texture[36][70] = 1;	doodle_right_transparency_texture[36][71] = 1;	doodle_right_transparency_texture[36][72] = 1;	doodle_right_transparency_texture[36][73] = 1;	doodle_right_transparency_texture[36][74] = 1;	doodle_right_transparency_texture[36][75] = 1;	doodle_right_transparency_texture[36][76] = 1;	doodle_right_transparency_texture[36][77] = 1;	doodle_right_transparency_texture[36][78] = 1;	doodle_right_transparency_texture[36][79] = 1;	doodle_right_transparency_texture[37][0] = 1;	doodle_right_transparency_texture[37][1] = 1;	doodle_right_transparency_texture[37][2] = 1;	doodle_right_transparency_texture[37][3] = 1;	doodle_right_transparency_texture[37][4] = 0;	doodle_right_transparency_texture[37][5] = 0;	doodle_right_transparency_texture[37][6] = 0;	doodle_right_transparency_texture[37][7] = 0;	doodle_right_transparency_texture[37][8] = 0;	doodle_right_transparency_texture[37][9] = 0;	doodle_right_transparency_texture[37][10] = 0;	doodle_right_transparency_texture[37][11] = 0;	doodle_right_transparency_texture[37][12] = 0;	doodle_right_transparency_texture[37][13] = 0;	doodle_right_transparency_texture[37][14] = 0;	doodle_right_transparency_texture[37][15] = 0;	doodle_right_transparency_texture[37][16] = 0;	doodle_right_transparency_texture[37][17] = 0;	doodle_right_transparency_texture[37][18] = 0;	doodle_right_transparency_texture[37][19] = 0;	doodle_right_transparency_texture[37][20] = 0;	doodle_right_transparency_texture[37][21] = 0;	doodle_right_transparency_texture[37][22] = 0;	doodle_right_transparency_texture[37][23] = 0;	doodle_right_transparency_texture[37][24] = 0;	doodle_right_transparency_texture[37][25] = 0;	doodle_right_transparency_texture[37][26] = 0;	doodle_right_transparency_texture[37][27] = 0;	doodle_right_transparency_texture[37][28] = 0;	doodle_right_transparency_texture[37][29] = 0;	doodle_right_transparency_texture[37][30] = 0;	doodle_right_transparency_texture[37][31] = 0;	doodle_right_transparency_texture[37][32] = 0;	doodle_right_transparency_texture[37][33] = 0;	doodle_right_transparency_texture[37][34] = 0;	doodle_right_transparency_texture[37][35] = 0;	doodle_right_transparency_texture[37][36] = 0;	doodle_right_transparency_texture[37][37] = 0;	doodle_right_transparency_texture[37][38] = 0;	doodle_right_transparency_texture[37][39] = 0;	doodle_right_transparency_texture[37][40] = 0;	doodle_right_transparency_texture[37][41] = 0;	doodle_right_transparency_texture[37][42] = 0;	doodle_right_transparency_texture[37][43] = 0;	doodle_right_transparency_texture[37][44] = 0;	doodle_right_transparency_texture[37][45] = 0;	doodle_right_transparency_texture[37][46] = 0;	doodle_right_transparency_texture[37][47] = 0;	doodle_right_transparency_texture[37][48] = 0;	doodle_right_transparency_texture[37][49] = 0;	doodle_right_transparency_texture[37][50] = 0;	doodle_right_transparency_texture[37][51] = 0;	doodle_right_transparency_texture[37][52] = 1;	doodle_right_transparency_texture[37][53] = 1;	doodle_right_transparency_texture[37][54] = 1;	doodle_right_transparency_texture[37][55] = 1;	doodle_right_transparency_texture[37][56] = 1;	doodle_right_transparency_texture[37][57] = 1;	doodle_right_transparency_texture[37][58] = 1;	doodle_right_transparency_texture[37][59] = 1;	doodle_right_transparency_texture[37][60] = 1;	doodle_right_transparency_texture[37][61] = 1;	doodle_right_transparency_texture[37][62] = 1;	doodle_right_transparency_texture[37][63] = 1;	doodle_right_transparency_texture[37][64] = 1;	doodle_right_transparency_texture[37][65] = 1;	doodle_right_transparency_texture[37][66] = 1;	doodle_right_transparency_texture[37][67] = 1;	doodle_right_transparency_texture[37][68] = 1;	doodle_right_transparency_texture[37][69] = 1;	doodle_right_transparency_texture[37][70] = 1;	doodle_right_transparency_texture[37][71] = 1;	doodle_right_transparency_texture[37][72] = 1;	doodle_right_transparency_texture[37][73] = 1;	doodle_right_transparency_texture[37][74] = 1;	doodle_right_transparency_texture[37][75] = 1;	doodle_right_transparency_texture[37][76] = 1;	doodle_right_transparency_texture[37][77] = 1;	doodle_right_transparency_texture[37][78] = 1;	doodle_right_transparency_texture[37][79] = 1;	doodle_right_transparency_texture[38][0] = 1;	doodle_right_transparency_texture[38][1] = 1;	doodle_right_transparency_texture[38][2] = 1;	doodle_right_transparency_texture[38][3] = 1;	doodle_right_transparency_texture[38][4] = 0;	doodle_right_transparency_texture[38][5] = 0;	doodle_right_transparency_texture[38][6] = 0;	doodle_right_transparency_texture[38][7] = 0;	doodle_right_transparency_texture[38][8] = 0;	doodle_right_transparency_texture[38][9] = 0;	doodle_right_transparency_texture[38][10] = 0;	doodle_right_transparency_texture[38][11] = 0;	doodle_right_transparency_texture[38][12] = 0;	doodle_right_transparency_texture[38][13] = 0;	doodle_right_transparency_texture[38][14] = 0;	doodle_right_transparency_texture[38][15] = 0;	doodle_right_transparency_texture[38][16] = 0;	doodle_right_transparency_texture[38][17] = 0;	doodle_right_transparency_texture[38][18] = 0;	doodle_right_transparency_texture[38][19] = 0;	doodle_right_transparency_texture[38][20] = 0;	doodle_right_transparency_texture[38][21] = 0;	doodle_right_transparency_texture[38][22] = 0;	doodle_right_transparency_texture[38][23] = 0;	doodle_right_transparency_texture[38][24] = 0;	doodle_right_transparency_texture[38][25] = 0;	doodle_right_transparency_texture[38][26] = 0;	doodle_right_transparency_texture[38][27] = 0;	doodle_right_transparency_texture[38][28] = 0;	doodle_right_transparency_texture[38][29] = 0;	doodle_right_transparency_texture[38][30] = 0;	doodle_right_transparency_texture[38][31] = 0;	doodle_right_transparency_texture[38][32] = 0;	doodle_right_transparency_texture[38][33] = 0;	doodle_right_transparency_texture[38][34] = 0;	doodle_right_transparency_texture[38][35] = 0;	doodle_right_transparency_texture[38][36] = 0;	doodle_right_transparency_texture[38][37] = 0;	doodle_right_transparency_texture[38][38] = 0;	doodle_right_transparency_texture[38][39] = 0;	doodle_right_transparency_texture[38][40] = 0;	doodle_right_transparency_texture[38][41] = 0;	doodle_right_transparency_texture[38][42] = 0;	doodle_right_transparency_texture[38][43] = 0;	doodle_right_transparency_texture[38][44] = 0;	doodle_right_transparency_texture[38][45] = 0;	doodle_right_transparency_texture[38][46] = 0;	doodle_right_transparency_texture[38][47] = 0;	doodle_right_transparency_texture[38][48] = 0;	doodle_right_transparency_texture[38][49] = 0;	doodle_right_transparency_texture[38][50] = 0;	doodle_right_transparency_texture[38][51] = 0;	doodle_right_transparency_texture[38][52] = 1;	doodle_right_transparency_texture[38][53] = 1;	doodle_right_transparency_texture[38][54] = 1;	doodle_right_transparency_texture[38][55] = 1;	doodle_right_transparency_texture[38][56] = 1;	doodle_right_transparency_texture[38][57] = 1;	doodle_right_transparency_texture[38][58] = 1;	doodle_right_transparency_texture[38][59] = 1;	doodle_right_transparency_texture[38][60] = 1;	doodle_right_transparency_texture[38][61] = 1;	doodle_right_transparency_texture[38][62] = 1;	doodle_right_transparency_texture[38][63] = 1;	doodle_right_transparency_texture[38][64] = 1;	doodle_right_transparency_texture[38][65] = 1;	doodle_right_transparency_texture[38][66] = 1;	doodle_right_transparency_texture[38][67] = 1;	doodle_right_transparency_texture[38][68] = 1;	doodle_right_transparency_texture[38][69] = 1;	doodle_right_transparency_texture[38][70] = 1;	doodle_right_transparency_texture[38][71] = 1;	doodle_right_transparency_texture[38][72] = 1;	doodle_right_transparency_texture[38][73] = 1;	doodle_right_transparency_texture[38][74] = 1;	doodle_right_transparency_texture[38][75] = 1;	doodle_right_transparency_texture[38][76] = 1;	doodle_right_transparency_texture[38][77] = 1;	doodle_right_transparency_texture[38][78] = 1;	doodle_right_transparency_texture[38][79] = 1;	doodle_right_transparency_texture[39][0] = 1;	doodle_right_transparency_texture[39][1] = 1;	doodle_right_transparency_texture[39][2] = 1;	doodle_right_transparency_texture[39][3] = 1;	doodle_right_transparency_texture[39][4] = 0;	doodle_right_transparency_texture[39][5] = 0;	doodle_right_transparency_texture[39][6] = 0;	doodle_right_transparency_texture[39][7] = 0;	doodle_right_transparency_texture[39][8] = 0;	doodle_right_transparency_texture[39][9] = 0;	doodle_right_transparency_texture[39][10] = 0;	doodle_right_transparency_texture[39][11] = 0;	doodle_right_transparency_texture[39][12] = 0;	doodle_right_transparency_texture[39][13] = 0;	doodle_right_transparency_texture[39][14] = 0;	doodle_right_transparency_texture[39][15] = 0;	doodle_right_transparency_texture[39][16] = 0;	doodle_right_transparency_texture[39][17] = 0;	doodle_right_transparency_texture[39][18] = 0;	doodle_right_transparency_texture[39][19] = 0;	doodle_right_transparency_texture[39][20] = 0;	doodle_right_transparency_texture[39][21] = 0;	doodle_right_transparency_texture[39][22] = 0;	doodle_right_transparency_texture[39][23] = 0;	doodle_right_transparency_texture[39][24] = 0;	doodle_right_transparency_texture[39][25] = 0;	doodle_right_transparency_texture[39][26] = 0;	doodle_right_transparency_texture[39][27] = 0;	doodle_right_transparency_texture[39][28] = 0;	doodle_right_transparency_texture[39][29] = 0;	doodle_right_transparency_texture[39][30] = 0;	doodle_right_transparency_texture[39][31] = 0;	doodle_right_transparency_texture[39][32] = 0;	doodle_right_transparency_texture[39][33] = 0;	doodle_right_transparency_texture[39][34] = 0;	doodle_right_transparency_texture[39][35] = 0;	doodle_right_transparency_texture[39][36] = 0;	doodle_right_transparency_texture[39][37] = 0;	doodle_right_transparency_texture[39][38] = 0;	doodle_right_transparency_texture[39][39] = 0;	doodle_right_transparency_texture[39][40] = 0;	doodle_right_transparency_texture[39][41] = 0;	doodle_right_transparency_texture[39][42] = 0;	doodle_right_transparency_texture[39][43] = 0;	doodle_right_transparency_texture[39][44] = 0;	doodle_right_transparency_texture[39][45] = 0;	doodle_right_transparency_texture[39][46] = 0;	doodle_right_transparency_texture[39][47] = 0;	doodle_right_transparency_texture[39][48] = 0;	doodle_right_transparency_texture[39][49] = 0;	doodle_right_transparency_texture[39][50] = 0;	doodle_right_transparency_texture[39][51] = 0;	doodle_right_transparency_texture[39][52] = 1;	doodle_right_transparency_texture[39][53] = 1;	doodle_right_transparency_texture[39][54] = 1;	doodle_right_transparency_texture[39][55] = 1;	doodle_right_transparency_texture[39][56] = 1;	doodle_right_transparency_texture[39][57] = 1;	doodle_right_transparency_texture[39][58] = 1;	doodle_right_transparency_texture[39][59] = 1;	doodle_right_transparency_texture[39][60] = 1;	doodle_right_transparency_texture[39][61] = 1;	doodle_right_transparency_texture[39][62] = 1;	doodle_right_transparency_texture[39][63] = 1;	doodle_right_transparency_texture[39][64] = 1;	doodle_right_transparency_texture[39][65] = 1;	doodle_right_transparency_texture[39][66] = 1;	doodle_right_transparency_texture[39][67] = 1;	doodle_right_transparency_texture[39][68] = 1;	doodle_right_transparency_texture[39][69] = 1;	doodle_right_transparency_texture[39][70] = 1;	doodle_right_transparency_texture[39][71] = 1;	doodle_right_transparency_texture[39][72] = 1;	doodle_right_transparency_texture[39][73] = 1;	doodle_right_transparency_texture[39][74] = 1;	doodle_right_transparency_texture[39][75] = 1;	doodle_right_transparency_texture[39][76] = 1;	doodle_right_transparency_texture[39][77] = 1;	doodle_right_transparency_texture[39][78] = 1;	doodle_right_transparency_texture[39][79] = 1;	doodle_right_transparency_texture[40][0] = 1;	doodle_right_transparency_texture[40][1] = 1;	doodle_right_transparency_texture[40][2] = 1;	doodle_right_transparency_texture[40][3] = 1;	doodle_right_transparency_texture[40][4] = 0;	doodle_right_transparency_texture[40][5] = 0;	doodle_right_transparency_texture[40][6] = 0;	doodle_right_transparency_texture[40][7] = 0;	doodle_right_transparency_texture[40][8] = 0;	doodle_right_transparency_texture[40][9] = 0;	doodle_right_transparency_texture[40][10] = 0;	doodle_right_transparency_texture[40][11] = 0;	doodle_right_transparency_texture[40][12] = 0;	doodle_right_transparency_texture[40][13] = 0;	doodle_right_transparency_texture[40][14] = 0;	doodle_right_transparency_texture[40][15] = 0;	doodle_right_transparency_texture[40][16] = 0;	doodle_right_transparency_texture[40][17] = 0;	doodle_right_transparency_texture[40][18] = 0;	doodle_right_transparency_texture[40][19] = 0;	doodle_right_transparency_texture[40][20] = 0;	doodle_right_transparency_texture[40][21] = 0;	doodle_right_transparency_texture[40][22] = 0;	doodle_right_transparency_texture[40][23] = 0;	doodle_right_transparency_texture[40][24] = 0;	doodle_right_transparency_texture[40][25] = 0;	doodle_right_transparency_texture[40][26] = 0;	doodle_right_transparency_texture[40][27] = 0;	doodle_right_transparency_texture[40][28] = 0;	doodle_right_transparency_texture[40][29] = 0;	doodle_right_transparency_texture[40][30] = 0;	doodle_right_transparency_texture[40][31] = 0;	doodle_right_transparency_texture[40][32] = 0;	doodle_right_transparency_texture[40][33] = 0;	doodle_right_transparency_texture[40][34] = 0;	doodle_right_transparency_texture[40][35] = 0;	doodle_right_transparency_texture[40][36] = 0;	doodle_right_transparency_texture[40][37] = 0;	doodle_right_transparency_texture[40][38] = 0;	doodle_right_transparency_texture[40][39] = 0;	doodle_right_transparency_texture[40][40] = 0;	doodle_right_transparency_texture[40][41] = 0;	doodle_right_transparency_texture[40][42] = 0;	doodle_right_transparency_texture[40][43] = 0;	doodle_right_transparency_texture[40][44] = 0;	doodle_right_transparency_texture[40][45] = 0;	doodle_right_transparency_texture[40][46] = 0;	doodle_right_transparency_texture[40][47] = 0;	doodle_right_transparency_texture[40][48] = 0;	doodle_right_transparency_texture[40][49] = 0;	doodle_right_transparency_texture[40][50] = 0;	doodle_right_transparency_texture[40][51] = 0;	doodle_right_transparency_texture[40][52] = 1;	doodle_right_transparency_texture[40][53] = 1;	doodle_right_transparency_texture[40][54] = 1;	doodle_right_transparency_texture[40][55] = 1;	doodle_right_transparency_texture[40][56] = 1;	doodle_right_transparency_texture[40][57] = 1;	doodle_right_transparency_texture[40][58] = 1;	doodle_right_transparency_texture[40][59] = 1;	doodle_right_transparency_texture[40][60] = 1;	doodle_right_transparency_texture[40][61] = 1;	doodle_right_transparency_texture[40][62] = 1;	doodle_right_transparency_texture[40][63] = 1;	doodle_right_transparency_texture[40][64] = 1;	doodle_right_transparency_texture[40][65] = 1;	doodle_right_transparency_texture[40][66] = 1;	doodle_right_transparency_texture[40][67] = 1;	doodle_right_transparency_texture[40][68] = 1;	doodle_right_transparency_texture[40][69] = 1;	doodle_right_transparency_texture[40][70] = 1;	doodle_right_transparency_texture[40][71] = 1;	doodle_right_transparency_texture[40][72] = 1;	doodle_right_transparency_texture[40][73] = 1;	doodle_right_transparency_texture[40][74] = 1;	doodle_right_transparency_texture[40][75] = 1;	doodle_right_transparency_texture[40][76] = 1;	doodle_right_transparency_texture[40][77] = 1;	doodle_right_transparency_texture[40][78] = 1;	doodle_right_transparency_texture[40][79] = 1;	doodle_right_transparency_texture[41][0] = 1;	doodle_right_transparency_texture[41][1] = 1;	doodle_right_transparency_texture[41][2] = 1;	doodle_right_transparency_texture[41][3] = 1;	doodle_right_transparency_texture[41][4] = 0;	doodle_right_transparency_texture[41][5] = 0;	doodle_right_transparency_texture[41][6] = 0;	doodle_right_transparency_texture[41][7] = 0;	doodle_right_transparency_texture[41][8] = 0;	doodle_right_transparency_texture[41][9] = 0;	doodle_right_transparency_texture[41][10] = 0;	doodle_right_transparency_texture[41][11] = 0;	doodle_right_transparency_texture[41][12] = 0;	doodle_right_transparency_texture[41][13] = 0;	doodle_right_transparency_texture[41][14] = 0;	doodle_right_transparency_texture[41][15] = 0;	doodle_right_transparency_texture[41][16] = 0;	doodle_right_transparency_texture[41][17] = 0;	doodle_right_transparency_texture[41][18] = 0;	doodle_right_transparency_texture[41][19] = 0;	doodle_right_transparency_texture[41][20] = 0;	doodle_right_transparency_texture[41][21] = 0;	doodle_right_transparency_texture[41][22] = 0;	doodle_right_transparency_texture[41][23] = 0;	doodle_right_transparency_texture[41][24] = 0;	doodle_right_transparency_texture[41][25] = 0;	doodle_right_transparency_texture[41][26] = 0;	doodle_right_transparency_texture[41][27] = 0;	doodle_right_transparency_texture[41][28] = 0;	doodle_right_transparency_texture[41][29] = 0;	doodle_right_transparency_texture[41][30] = 0;	doodle_right_transparency_texture[41][31] = 0;	doodle_right_transparency_texture[41][32] = 0;	doodle_right_transparency_texture[41][33] = 0;	doodle_right_transparency_texture[41][34] = 0;	doodle_right_transparency_texture[41][35] = 0;	doodle_right_transparency_texture[41][36] = 0;	doodle_right_transparency_texture[41][37] = 0;	doodle_right_transparency_texture[41][38] = 0;	doodle_right_transparency_texture[41][39] = 0;	doodle_right_transparency_texture[41][40] = 0;	doodle_right_transparency_texture[41][41] = 0;	doodle_right_transparency_texture[41][42] = 0;	doodle_right_transparency_texture[41][43] = 0;	doodle_right_transparency_texture[41][44] = 0;	doodle_right_transparency_texture[41][45] = 0;	doodle_right_transparency_texture[41][46] = 0;	doodle_right_transparency_texture[41][47] = 0;	doodle_right_transparency_texture[41][48] = 0;	doodle_right_transparency_texture[41][49] = 0;	doodle_right_transparency_texture[41][50] = 0;	doodle_right_transparency_texture[41][51] = 0;	doodle_right_transparency_texture[41][52] = 1;	doodle_right_transparency_texture[41][53] = 1;	doodle_right_transparency_texture[41][54] = 1;	doodle_right_transparency_texture[41][55] = 1;	doodle_right_transparency_texture[41][56] = 1;	doodle_right_transparency_texture[41][57] = 1;	doodle_right_transparency_texture[41][58] = 1;	doodle_right_transparency_texture[41][59] = 1;	doodle_right_transparency_texture[41][60] = 1;	doodle_right_transparency_texture[41][61] = 1;	doodle_right_transparency_texture[41][62] = 1;	doodle_right_transparency_texture[41][63] = 1;	doodle_right_transparency_texture[41][64] = 1;	doodle_right_transparency_texture[41][65] = 1;	doodle_right_transparency_texture[41][66] = 1;	doodle_right_transparency_texture[41][67] = 1;	doodle_right_transparency_texture[41][68] = 1;	doodle_right_transparency_texture[41][69] = 1;	doodle_right_transparency_texture[41][70] = 1;	doodle_right_transparency_texture[41][71] = 1;	doodle_right_transparency_texture[41][72] = 1;	doodle_right_transparency_texture[41][73] = 1;	doodle_right_transparency_texture[41][74] = 1;	doodle_right_transparency_texture[41][75] = 1;	doodle_right_transparency_texture[41][76] = 1;	doodle_right_transparency_texture[41][77] = 1;	doodle_right_transparency_texture[41][78] = 1;	doodle_right_transparency_texture[41][79] = 1;	doodle_right_transparency_texture[42][0] = 1;	doodle_right_transparency_texture[42][1] = 1;	doodle_right_transparency_texture[42][2] = 1;	doodle_right_transparency_texture[42][3] = 1;	doodle_right_transparency_texture[42][4] = 0;	doodle_right_transparency_texture[42][5] = 0;	doodle_right_transparency_texture[42][6] = 0;	doodle_right_transparency_texture[42][7] = 0;	doodle_right_transparency_texture[42][8] = 0;	doodle_right_transparency_texture[42][9] = 0;	doodle_right_transparency_texture[42][10] = 0;	doodle_right_transparency_texture[42][11] = 0;	doodle_right_transparency_texture[42][12] = 0;	doodle_right_transparency_texture[42][13] = 0;	doodle_right_transparency_texture[42][14] = 0;	doodle_right_transparency_texture[42][15] = 0;	doodle_right_transparency_texture[42][16] = 0;	doodle_right_transparency_texture[42][17] = 0;	doodle_right_transparency_texture[42][18] = 0;	doodle_right_transparency_texture[42][19] = 0;	doodle_right_transparency_texture[42][20] = 0;	doodle_right_transparency_texture[42][21] = 0;	doodle_right_transparency_texture[42][22] = 0;	doodle_right_transparency_texture[42][23] = 0;	doodle_right_transparency_texture[42][24] = 0;	doodle_right_transparency_texture[42][25] = 0;	doodle_right_transparency_texture[42][26] = 0;	doodle_right_transparency_texture[42][27] = 0;	doodle_right_transparency_texture[42][28] = 0;	doodle_right_transparency_texture[42][29] = 0;	doodle_right_transparency_texture[42][30] = 0;	doodle_right_transparency_texture[42][31] = 0;	doodle_right_transparency_texture[42][32] = 0;	doodle_right_transparency_texture[42][33] = 0;	doodle_right_transparency_texture[42][34] = 0;	doodle_right_transparency_texture[42][35] = 0;	doodle_right_transparency_texture[42][36] = 0;	doodle_right_transparency_texture[42][37] = 0;	doodle_right_transparency_texture[42][38] = 0;	doodle_right_transparency_texture[42][39] = 0;	doodle_right_transparency_texture[42][40] = 0;	doodle_right_transparency_texture[42][41] = 0;	doodle_right_transparency_texture[42][42] = 0;	doodle_right_transparency_texture[42][43] = 0;	doodle_right_transparency_texture[42][44] = 0;	doodle_right_transparency_texture[42][45] = 0;	doodle_right_transparency_texture[42][46] = 0;	doodle_right_transparency_texture[42][47] = 0;	doodle_right_transparency_texture[42][48] = 0;	doodle_right_transparency_texture[42][49] = 0;	doodle_right_transparency_texture[42][50] = 0;	doodle_right_transparency_texture[42][51] = 0;	doodle_right_transparency_texture[42][52] = 1;	doodle_right_transparency_texture[42][53] = 1;	doodle_right_transparency_texture[42][54] = 1;	doodle_right_transparency_texture[42][55] = 1;	doodle_right_transparency_texture[42][56] = 1;	doodle_right_transparency_texture[42][57] = 1;	doodle_right_transparency_texture[42][58] = 1;	doodle_right_transparency_texture[42][59] = 1;	doodle_right_transparency_texture[42][60] = 1;	doodle_right_transparency_texture[42][61] = 1;	doodle_right_transparency_texture[42][62] = 1;	doodle_right_transparency_texture[42][63] = 1;	doodle_right_transparency_texture[42][64] = 1;	doodle_right_transparency_texture[42][65] = 1;	doodle_right_transparency_texture[42][66] = 1;	doodle_right_transparency_texture[42][67] = 1;	doodle_right_transparency_texture[42][68] = 1;	doodle_right_transparency_texture[42][69] = 1;	doodle_right_transparency_texture[42][70] = 1;	doodle_right_transparency_texture[42][71] = 1;	doodle_right_transparency_texture[42][72] = 1;	doodle_right_transparency_texture[42][73] = 1;	doodle_right_transparency_texture[42][74] = 1;	doodle_right_transparency_texture[42][75] = 1;	doodle_right_transparency_texture[42][76] = 1;	doodle_right_transparency_texture[42][77] = 1;	doodle_right_transparency_texture[42][78] = 1;	doodle_right_transparency_texture[42][79] = 1;	doodle_right_transparency_texture[43][0] = 1;	doodle_right_transparency_texture[43][1] = 1;	doodle_right_transparency_texture[43][2] = 1;	doodle_right_transparency_texture[43][3] = 1;	doodle_right_transparency_texture[43][4] = 0;	doodle_right_transparency_texture[43][5] = 0;	doodle_right_transparency_texture[43][6] = 0;	doodle_right_transparency_texture[43][7] = 0;	doodle_right_transparency_texture[43][8] = 0;	doodle_right_transparency_texture[43][9] = 0;	doodle_right_transparency_texture[43][10] = 0;	doodle_right_transparency_texture[43][11] = 0;	doodle_right_transparency_texture[43][12] = 0;	doodle_right_transparency_texture[43][13] = 0;	doodle_right_transparency_texture[43][14] = 0;	doodle_right_transparency_texture[43][15] = 0;	doodle_right_transparency_texture[43][16] = 0;	doodle_right_transparency_texture[43][17] = 0;	doodle_right_transparency_texture[43][18] = 0;	doodle_right_transparency_texture[43][19] = 0;	doodle_right_transparency_texture[43][20] = 0;	doodle_right_transparency_texture[43][21] = 0;	doodle_right_transparency_texture[43][22] = 0;	doodle_right_transparency_texture[43][23] = 0;	doodle_right_transparency_texture[43][24] = 0;	doodle_right_transparency_texture[43][25] = 0;	doodle_right_transparency_texture[43][26] = 0;	doodle_right_transparency_texture[43][27] = 0;	doodle_right_transparency_texture[43][28] = 0;	doodle_right_transparency_texture[43][29] = 0;	doodle_right_transparency_texture[43][30] = 0;	doodle_right_transparency_texture[43][31] = 0;	doodle_right_transparency_texture[43][32] = 0;	doodle_right_transparency_texture[43][33] = 0;	doodle_right_transparency_texture[43][34] = 0;	doodle_right_transparency_texture[43][35] = 0;	doodle_right_transparency_texture[43][36] = 0;	doodle_right_transparency_texture[43][37] = 0;	doodle_right_transparency_texture[43][38] = 0;	doodle_right_transparency_texture[43][39] = 0;	doodle_right_transparency_texture[43][40] = 0;	doodle_right_transparency_texture[43][41] = 0;	doodle_right_transparency_texture[43][42] = 0;	doodle_right_transparency_texture[43][43] = 0;	doodle_right_transparency_texture[43][44] = 0;	doodle_right_transparency_texture[43][45] = 0;	doodle_right_transparency_texture[43][46] = 0;	doodle_right_transparency_texture[43][47] = 0;	doodle_right_transparency_texture[43][48] = 0;	doodle_right_transparency_texture[43][49] = 0;	doodle_right_transparency_texture[43][50] = 0;	doodle_right_transparency_texture[43][51] = 0;	doodle_right_transparency_texture[43][52] = 1;	doodle_right_transparency_texture[43][53] = 1;	doodle_right_transparency_texture[43][54] = 1;	doodle_right_transparency_texture[43][55] = 1;	doodle_right_transparency_texture[43][56] = 1;	doodle_right_transparency_texture[43][57] = 1;	doodle_right_transparency_texture[43][58] = 1;	doodle_right_transparency_texture[43][59] = 1;	doodle_right_transparency_texture[43][60] = 1;	doodle_right_transparency_texture[43][61] = 1;	doodle_right_transparency_texture[43][62] = 1;	doodle_right_transparency_texture[43][63] = 1;	doodle_right_transparency_texture[43][64] = 1;	doodle_right_transparency_texture[43][65] = 1;	doodle_right_transparency_texture[43][66] = 1;	doodle_right_transparency_texture[43][67] = 1;	doodle_right_transparency_texture[43][68] = 1;	doodle_right_transparency_texture[43][69] = 1;	doodle_right_transparency_texture[43][70] = 1;	doodle_right_transparency_texture[43][71] = 1;	doodle_right_transparency_texture[43][72] = 1;	doodle_right_transparency_texture[43][73] = 1;	doodle_right_transparency_texture[43][74] = 1;	doodle_right_transparency_texture[43][75] = 1;	doodle_right_transparency_texture[43][76] = 1;	doodle_right_transparency_texture[43][77] = 1;	doodle_right_transparency_texture[43][78] = 1;	doodle_right_transparency_texture[43][79] = 1;	doodle_right_transparency_texture[44][0] = 1;	doodle_right_transparency_texture[44][1] = 1;	doodle_right_transparency_texture[44][2] = 1;	doodle_right_transparency_texture[44][3] = 1;	doodle_right_transparency_texture[44][4] = 0;	doodle_right_transparency_texture[44][5] = 0;	doodle_right_transparency_texture[44][6] = 0;	doodle_right_transparency_texture[44][7] = 0;	doodle_right_transparency_texture[44][8] = 0;	doodle_right_transparency_texture[44][9] = 0;	doodle_right_transparency_texture[44][10] = 0;	doodle_right_transparency_texture[44][11] = 0;	doodle_right_transparency_texture[44][12] = 0;	doodle_right_transparency_texture[44][13] = 0;	doodle_right_transparency_texture[44][14] = 0;	doodle_right_transparency_texture[44][15] = 0;	doodle_right_transparency_texture[44][16] = 0;	doodle_right_transparency_texture[44][17] = 0;	doodle_right_transparency_texture[44][18] = 0;	doodle_right_transparency_texture[44][19] = 0;	doodle_right_transparency_texture[44][20] = 0;	doodle_right_transparency_texture[44][21] = 0;	doodle_right_transparency_texture[44][22] = 0;	doodle_right_transparency_texture[44][23] = 0;	doodle_right_transparency_texture[44][24] = 0;	doodle_right_transparency_texture[44][25] = 0;	doodle_right_transparency_texture[44][26] = 0;	doodle_right_transparency_texture[44][27] = 0;	doodle_right_transparency_texture[44][28] = 0;	doodle_right_transparency_texture[44][29] = 0;	doodle_right_transparency_texture[44][30] = 0;	doodle_right_transparency_texture[44][31] = 0;	doodle_right_transparency_texture[44][32] = 0;	doodle_right_transparency_texture[44][33] = 0;	doodle_right_transparency_texture[44][34] = 0;	doodle_right_transparency_texture[44][35] = 0;	doodle_right_transparency_texture[44][36] = 0;	doodle_right_transparency_texture[44][37] = 0;	doodle_right_transparency_texture[44][38] = 0;	doodle_right_transparency_texture[44][39] = 0;	doodle_right_transparency_texture[44][40] = 0;	doodle_right_transparency_texture[44][41] = 0;	doodle_right_transparency_texture[44][42] = 0;	doodle_right_transparency_texture[44][43] = 0;	doodle_right_transparency_texture[44][44] = 0;	doodle_right_transparency_texture[44][45] = 0;	doodle_right_transparency_texture[44][46] = 0;	doodle_right_transparency_texture[44][47] = 0;	doodle_right_transparency_texture[44][48] = 0;	doodle_right_transparency_texture[44][49] = 0;	doodle_right_transparency_texture[44][50] = 0;	doodle_right_transparency_texture[44][51] = 0;	doodle_right_transparency_texture[44][52] = 1;	doodle_right_transparency_texture[44][53] = 1;	doodle_right_transparency_texture[44][54] = 1;	doodle_right_transparency_texture[44][55] = 1;	doodle_right_transparency_texture[44][56] = 1;	doodle_right_transparency_texture[44][57] = 1;	doodle_right_transparency_texture[44][58] = 1;	doodle_right_transparency_texture[44][59] = 1;	doodle_right_transparency_texture[44][60] = 1;	doodle_right_transparency_texture[44][61] = 1;	doodle_right_transparency_texture[44][62] = 1;	doodle_right_transparency_texture[44][63] = 1;	doodle_right_transparency_texture[44][64] = 1;	doodle_right_transparency_texture[44][65] = 1;	doodle_right_transparency_texture[44][66] = 1;	doodle_right_transparency_texture[44][67] = 1;	doodle_right_transparency_texture[44][68] = 1;	doodle_right_transparency_texture[44][69] = 1;	doodle_right_transparency_texture[44][70] = 1;	doodle_right_transparency_texture[44][71] = 1;	doodle_right_transparency_texture[44][72] = 1;	doodle_right_transparency_texture[44][73] = 1;	doodle_right_transparency_texture[44][74] = 1;	doodle_right_transparency_texture[44][75] = 1;	doodle_right_transparency_texture[44][76] = 1;	doodle_right_transparency_texture[44][77] = 1;	doodle_right_transparency_texture[44][78] = 1;	doodle_right_transparency_texture[44][79] = 1;	doodle_right_transparency_texture[45][0] = 1;	doodle_right_transparency_texture[45][1] = 1;	doodle_right_transparency_texture[45][2] = 1;	doodle_right_transparency_texture[45][3] = 1;	doodle_right_transparency_texture[45][4] = 0;	doodle_right_transparency_texture[45][5] = 0;	doodle_right_transparency_texture[45][6] = 0;	doodle_right_transparency_texture[45][7] = 0;	doodle_right_transparency_texture[45][8] = 0;	doodle_right_transparency_texture[45][9] = 0;	doodle_right_transparency_texture[45][10] = 0;	doodle_right_transparency_texture[45][11] = 0;	doodle_right_transparency_texture[45][12] = 0;	doodle_right_transparency_texture[45][13] = 0;	doodle_right_transparency_texture[45][14] = 0;	doodle_right_transparency_texture[45][15] = 0;	doodle_right_transparency_texture[45][16] = 0;	doodle_right_transparency_texture[45][17] = 0;	doodle_right_transparency_texture[45][18] = 0;	doodle_right_transparency_texture[45][19] = 0;	doodle_right_transparency_texture[45][20] = 0;	doodle_right_transparency_texture[45][21] = 0;	doodle_right_transparency_texture[45][22] = 0;	doodle_right_transparency_texture[45][23] = 0;	doodle_right_transparency_texture[45][24] = 0;	doodle_right_transparency_texture[45][25] = 0;	doodle_right_transparency_texture[45][26] = 0;	doodle_right_transparency_texture[45][27] = 0;	doodle_right_transparency_texture[45][28] = 0;	doodle_right_transparency_texture[45][29] = 0;	doodle_right_transparency_texture[45][30] = 0;	doodle_right_transparency_texture[45][31] = 0;	doodle_right_transparency_texture[45][32] = 0;	doodle_right_transparency_texture[45][33] = 0;	doodle_right_transparency_texture[45][34] = 0;	doodle_right_transparency_texture[45][35] = 0;	doodle_right_transparency_texture[45][36] = 0;	doodle_right_transparency_texture[45][37] = 0;	doodle_right_transparency_texture[45][38] = 0;	doodle_right_transparency_texture[45][39] = 0;	doodle_right_transparency_texture[45][40] = 0;	doodle_right_transparency_texture[45][41] = 0;	doodle_right_transparency_texture[45][42] = 0;	doodle_right_transparency_texture[45][43] = 0;	doodle_right_transparency_texture[45][44] = 0;	doodle_right_transparency_texture[45][45] = 0;	doodle_right_transparency_texture[45][46] = 0;	doodle_right_transparency_texture[45][47] = 0;	doodle_right_transparency_texture[45][48] = 0;	doodle_right_transparency_texture[45][49] = 0;	doodle_right_transparency_texture[45][50] = 0;	doodle_right_transparency_texture[45][51] = 0;	doodle_right_transparency_texture[45][52] = 1;	doodle_right_transparency_texture[45][53] = 1;	doodle_right_transparency_texture[45][54] = 1;	doodle_right_transparency_texture[45][55] = 1;	doodle_right_transparency_texture[45][56] = 1;	doodle_right_transparency_texture[45][57] = 1;	doodle_right_transparency_texture[45][58] = 1;	doodle_right_transparency_texture[45][59] = 1;	doodle_right_transparency_texture[45][60] = 1;	doodle_right_transparency_texture[45][61] = 1;	doodle_right_transparency_texture[45][62] = 1;	doodle_right_transparency_texture[45][63] = 1;	doodle_right_transparency_texture[45][64] = 1;	doodle_right_transparency_texture[45][65] = 1;	doodle_right_transparency_texture[45][66] = 1;	doodle_right_transparency_texture[45][67] = 1;	doodle_right_transparency_texture[45][68] = 1;	doodle_right_transparency_texture[45][69] = 1;	doodle_right_transparency_texture[45][70] = 1;	doodle_right_transparency_texture[45][71] = 1;	doodle_right_transparency_texture[45][72] = 1;	doodle_right_transparency_texture[45][73] = 1;	doodle_right_transparency_texture[45][74] = 1;	doodle_right_transparency_texture[45][75] = 1;	doodle_right_transparency_texture[45][76] = 1;	doodle_right_transparency_texture[45][77] = 1;	doodle_right_transparency_texture[45][78] = 1;	doodle_right_transparency_texture[45][79] = 1;	doodle_right_transparency_texture[46][0] = 1;	doodle_right_transparency_texture[46][1] = 1;	doodle_right_transparency_texture[46][2] = 1;	doodle_right_transparency_texture[46][3] = 1;	doodle_right_transparency_texture[46][4] = 0;	doodle_right_transparency_texture[46][5] = 0;	doodle_right_transparency_texture[46][6] = 0;	doodle_right_transparency_texture[46][7] = 0;	doodle_right_transparency_texture[46][8] = 0;	doodle_right_transparency_texture[46][9] = 0;	doodle_right_transparency_texture[46][10] = 0;	doodle_right_transparency_texture[46][11] = 0;	doodle_right_transparency_texture[46][12] = 0;	doodle_right_transparency_texture[46][13] = 0;	doodle_right_transparency_texture[46][14] = 0;	doodle_right_transparency_texture[46][15] = 0;	doodle_right_transparency_texture[46][16] = 0;	doodle_right_transparency_texture[46][17] = 0;	doodle_right_transparency_texture[46][18] = 0;	doodle_right_transparency_texture[46][19] = 0;	doodle_right_transparency_texture[46][20] = 0;	doodle_right_transparency_texture[46][21] = 0;	doodle_right_transparency_texture[46][22] = 0;	doodle_right_transparency_texture[46][23] = 0;	doodle_right_transparency_texture[46][24] = 0;	doodle_right_transparency_texture[46][25] = 0;	doodle_right_transparency_texture[46][26] = 0;	doodle_right_transparency_texture[46][27] = 0;	doodle_right_transparency_texture[46][28] = 0;	doodle_right_transparency_texture[46][29] = 0;	doodle_right_transparency_texture[46][30] = 0;	doodle_right_transparency_texture[46][31] = 0;	doodle_right_transparency_texture[46][32] = 0;	doodle_right_transparency_texture[46][33] = 0;	doodle_right_transparency_texture[46][34] = 0;	doodle_right_transparency_texture[46][35] = 0;	doodle_right_transparency_texture[46][36] = 0;	doodle_right_transparency_texture[46][37] = 0;	doodle_right_transparency_texture[46][38] = 0;	doodle_right_transparency_texture[46][39] = 0;	doodle_right_transparency_texture[46][40] = 0;	doodle_right_transparency_texture[46][41] = 0;	doodle_right_transparency_texture[46][42] = 0;	doodle_right_transparency_texture[46][43] = 0;	doodle_right_transparency_texture[46][44] = 0;	doodle_right_transparency_texture[46][45] = 0;	doodle_right_transparency_texture[46][46] = 0;	doodle_right_transparency_texture[46][47] = 0;	doodle_right_transparency_texture[46][48] = 0;	doodle_right_transparency_texture[46][49] = 0;	doodle_right_transparency_texture[46][50] = 0;	doodle_right_transparency_texture[46][51] = 0;	doodle_right_transparency_texture[46][52] = 1;	doodle_right_transparency_texture[46][53] = 1;	doodle_right_transparency_texture[46][54] = 1;	doodle_right_transparency_texture[46][55] = 1;	doodle_right_transparency_texture[46][56] = 1;	doodle_right_transparency_texture[46][57] = 1;	doodle_right_transparency_texture[46][58] = 1;	doodle_right_transparency_texture[46][59] = 1;	doodle_right_transparency_texture[46][60] = 1;	doodle_right_transparency_texture[46][61] = 1;	doodle_right_transparency_texture[46][62] = 1;	doodle_right_transparency_texture[46][63] = 1;	doodle_right_transparency_texture[46][64] = 1;	doodle_right_transparency_texture[46][65] = 1;	doodle_right_transparency_texture[46][66] = 1;	doodle_right_transparency_texture[46][67] = 1;	doodle_right_transparency_texture[46][68] = 1;	doodle_right_transparency_texture[46][69] = 1;	doodle_right_transparency_texture[46][70] = 1;	doodle_right_transparency_texture[46][71] = 1;	doodle_right_transparency_texture[46][72] = 1;	doodle_right_transparency_texture[46][73] = 1;	doodle_right_transparency_texture[46][74] = 1;	doodle_right_transparency_texture[46][75] = 1;	doodle_right_transparency_texture[46][76] = 1;	doodle_right_transparency_texture[46][77] = 1;	doodle_right_transparency_texture[46][78] = 1;	doodle_right_transparency_texture[46][79] = 1;	doodle_right_transparency_texture[47][0] = 1;	doodle_right_transparency_texture[47][1] = 1;	doodle_right_transparency_texture[47][2] = 1;	doodle_right_transparency_texture[47][3] = 1;	doodle_right_transparency_texture[47][4] = 0;	doodle_right_transparency_texture[47][5] = 0;	doodle_right_transparency_texture[47][6] = 0;	doodle_right_transparency_texture[47][7] = 0;	doodle_right_transparency_texture[47][8] = 0;	doodle_right_transparency_texture[47][9] = 0;	doodle_right_transparency_texture[47][10] = 0;	doodle_right_transparency_texture[47][11] = 0;	doodle_right_transparency_texture[47][12] = 0;	doodle_right_transparency_texture[47][13] = 0;	doodle_right_transparency_texture[47][14] = 0;	doodle_right_transparency_texture[47][15] = 0;	doodle_right_transparency_texture[47][16] = 0;	doodle_right_transparency_texture[47][17] = 0;	doodle_right_transparency_texture[47][18] = 0;	doodle_right_transparency_texture[47][19] = 0;	doodle_right_transparency_texture[47][20] = 0;	doodle_right_transparency_texture[47][21] = 0;	doodle_right_transparency_texture[47][22] = 0;	doodle_right_transparency_texture[47][23] = 0;	doodle_right_transparency_texture[47][24] = 0;	doodle_right_transparency_texture[47][25] = 0;	doodle_right_transparency_texture[47][26] = 0;	doodle_right_transparency_texture[47][27] = 0;	doodle_right_transparency_texture[47][28] = 0;	doodle_right_transparency_texture[47][29] = 0;	doodle_right_transparency_texture[47][30] = 0;	doodle_right_transparency_texture[47][31] = 0;	doodle_right_transparency_texture[47][32] = 0;	doodle_right_transparency_texture[47][33] = 0;	doodle_right_transparency_texture[47][34] = 0;	doodle_right_transparency_texture[47][35] = 0;	doodle_right_transparency_texture[47][36] = 0;	doodle_right_transparency_texture[47][37] = 0;	doodle_right_transparency_texture[47][38] = 0;	doodle_right_transparency_texture[47][39] = 0;	doodle_right_transparency_texture[47][40] = 0;	doodle_right_transparency_texture[47][41] = 0;	doodle_right_transparency_texture[47][42] = 0;	doodle_right_transparency_texture[47][43] = 0;	doodle_right_transparency_texture[47][44] = 0;	doodle_right_transparency_texture[47][45] = 0;	doodle_right_transparency_texture[47][46] = 0;	doodle_right_transparency_texture[47][47] = 0;	doodle_right_transparency_texture[47][48] = 0;	doodle_right_transparency_texture[47][49] = 0;	doodle_right_transparency_texture[47][50] = 0;	doodle_right_transparency_texture[47][51] = 0;	doodle_right_transparency_texture[47][52] = 1;	doodle_right_transparency_texture[47][53] = 1;	doodle_right_transparency_texture[47][54] = 1;	doodle_right_transparency_texture[47][55] = 1;	doodle_right_transparency_texture[47][56] = 1;	doodle_right_transparency_texture[47][57] = 1;	doodle_right_transparency_texture[47][58] = 1;	doodle_right_transparency_texture[47][59] = 1;	doodle_right_transparency_texture[47][60] = 1;	doodle_right_transparency_texture[47][61] = 1;	doodle_right_transparency_texture[47][62] = 1;	doodle_right_transparency_texture[47][63] = 1;	doodle_right_transparency_texture[47][64] = 1;	doodle_right_transparency_texture[47][65] = 1;	doodle_right_transparency_texture[47][66] = 1;	doodle_right_transparency_texture[47][67] = 1;	doodle_right_transparency_texture[47][68] = 1;	doodle_right_transparency_texture[47][69] = 1;	doodle_right_transparency_texture[47][70] = 1;	doodle_right_transparency_texture[47][71] = 1;	doodle_right_transparency_texture[47][72] = 1;	doodle_right_transparency_texture[47][73] = 1;	doodle_right_transparency_texture[47][74] = 1;	doodle_right_transparency_texture[47][75] = 1;	doodle_right_transparency_texture[47][76] = 1;	doodle_right_transparency_texture[47][77] = 1;	doodle_right_transparency_texture[47][78] = 1;	doodle_right_transparency_texture[47][79] = 1;	doodle_right_transparency_texture[48][0] = 1;	doodle_right_transparency_texture[48][1] = 1;	doodle_right_transparency_texture[48][2] = 1;	doodle_right_transparency_texture[48][3] = 1;	doodle_right_transparency_texture[48][4] = 0;	doodle_right_transparency_texture[48][5] = 0;	doodle_right_transparency_texture[48][6] = 0;	doodle_right_transparency_texture[48][7] = 0;	doodle_right_transparency_texture[48][8] = 0;	doodle_right_transparency_texture[48][9] = 0;	doodle_right_transparency_texture[48][10] = 0;	doodle_right_transparency_texture[48][11] = 0;	doodle_right_transparency_texture[48][12] = 0;	doodle_right_transparency_texture[48][13] = 0;	doodle_right_transparency_texture[48][14] = 0;	doodle_right_transparency_texture[48][15] = 0;	doodle_right_transparency_texture[48][16] = 0;	doodle_right_transparency_texture[48][17] = 0;	doodle_right_transparency_texture[48][18] = 0;	doodle_right_transparency_texture[48][19] = 0;	doodle_right_transparency_texture[48][20] = 0;	doodle_right_transparency_texture[48][21] = 0;	doodle_right_transparency_texture[48][22] = 0;	doodle_right_transparency_texture[48][23] = 0;	doodle_right_transparency_texture[48][24] = 0;	doodle_right_transparency_texture[48][25] = 0;	doodle_right_transparency_texture[48][26] = 0;	doodle_right_transparency_texture[48][27] = 0;	doodle_right_transparency_texture[48][28] = 0;	doodle_right_transparency_texture[48][29] = 0;	doodle_right_transparency_texture[48][30] = 0;	doodle_right_transparency_texture[48][31] = 0;	doodle_right_transparency_texture[48][32] = 0;	doodle_right_transparency_texture[48][33] = 0;	doodle_right_transparency_texture[48][34] = 0;	doodle_right_transparency_texture[48][35] = 0;	doodle_right_transparency_texture[48][36] = 0;	doodle_right_transparency_texture[48][37] = 0;	doodle_right_transparency_texture[48][38] = 0;	doodle_right_transparency_texture[48][39] = 0;	doodle_right_transparency_texture[48][40] = 0;	doodle_right_transparency_texture[48][41] = 0;	doodle_right_transparency_texture[48][42] = 0;	doodle_right_transparency_texture[48][43] = 0;	doodle_right_transparency_texture[48][44] = 0;	doodle_right_transparency_texture[48][45] = 0;	doodle_right_transparency_texture[48][46] = 0;	doodle_right_transparency_texture[48][47] = 0;	doodle_right_transparency_texture[48][48] = 0;	doodle_right_transparency_texture[48][49] = 0;	doodle_right_transparency_texture[48][50] = 0;	doodle_right_transparency_texture[48][51] = 0;	doodle_right_transparency_texture[48][52] = 1;	doodle_right_transparency_texture[48][53] = 1;	doodle_right_transparency_texture[48][54] = 1;	doodle_right_transparency_texture[48][55] = 1;	doodle_right_transparency_texture[48][56] = 1;	doodle_right_transparency_texture[48][57] = 1;	doodle_right_transparency_texture[48][58] = 1;	doodle_right_transparency_texture[48][59] = 1;	doodle_right_transparency_texture[48][60] = 1;	doodle_right_transparency_texture[48][61] = 1;	doodle_right_transparency_texture[48][62] = 1;	doodle_right_transparency_texture[48][63] = 1;	doodle_right_transparency_texture[48][64] = 1;	doodle_right_transparency_texture[48][65] = 1;	doodle_right_transparency_texture[48][66] = 1;	doodle_right_transparency_texture[48][67] = 1;	doodle_right_transparency_texture[48][68] = 1;	doodle_right_transparency_texture[48][69] = 1;	doodle_right_transparency_texture[48][70] = 1;	doodle_right_transparency_texture[48][71] = 1;	doodle_right_transparency_texture[48][72] = 1;	doodle_right_transparency_texture[48][73] = 1;	doodle_right_transparency_texture[48][74] = 1;	doodle_right_transparency_texture[48][75] = 1;	doodle_right_transparency_texture[48][76] = 1;	doodle_right_transparency_texture[48][77] = 1;	doodle_right_transparency_texture[48][78] = 1;	doodle_right_transparency_texture[48][79] = 1;	doodle_right_transparency_texture[49][0] = 1;	doodle_right_transparency_texture[49][1] = 1;	doodle_right_transparency_texture[49][2] = 1;	doodle_right_transparency_texture[49][3] = 1;	doodle_right_transparency_texture[49][4] = 0;	doodle_right_transparency_texture[49][5] = 0;	doodle_right_transparency_texture[49][6] = 0;	doodle_right_transparency_texture[49][7] = 0;	doodle_right_transparency_texture[49][8] = 0;	doodle_right_transparency_texture[49][9] = 0;	doodle_right_transparency_texture[49][10] = 0;	doodle_right_transparency_texture[49][11] = 0;	doodle_right_transparency_texture[49][12] = 0;	doodle_right_transparency_texture[49][13] = 0;	doodle_right_transparency_texture[49][14] = 0;	doodle_right_transparency_texture[49][15] = 0;	doodle_right_transparency_texture[49][16] = 0;	doodle_right_transparency_texture[49][17] = 0;	doodle_right_transparency_texture[49][18] = 0;	doodle_right_transparency_texture[49][19] = 0;	doodle_right_transparency_texture[49][20] = 0;	doodle_right_transparency_texture[49][21] = 0;	doodle_right_transparency_texture[49][22] = 0;	doodle_right_transparency_texture[49][23] = 0;	doodle_right_transparency_texture[49][24] = 0;	doodle_right_transparency_texture[49][25] = 0;	doodle_right_transparency_texture[49][26] = 0;	doodle_right_transparency_texture[49][27] = 0;	doodle_right_transparency_texture[49][28] = 0;	doodle_right_transparency_texture[49][29] = 0;	doodle_right_transparency_texture[49][30] = 0;	doodle_right_transparency_texture[49][31] = 0;	doodle_right_transparency_texture[49][32] = 0;	doodle_right_transparency_texture[49][33] = 0;	doodle_right_transparency_texture[49][34] = 0;	doodle_right_transparency_texture[49][35] = 0;	doodle_right_transparency_texture[49][36] = 0;	doodle_right_transparency_texture[49][37] = 0;	doodle_right_transparency_texture[49][38] = 0;	doodle_right_transparency_texture[49][39] = 0;	doodle_right_transparency_texture[49][40] = 0;	doodle_right_transparency_texture[49][41] = 0;	doodle_right_transparency_texture[49][42] = 0;	doodle_right_transparency_texture[49][43] = 0;	doodle_right_transparency_texture[49][44] = 0;	doodle_right_transparency_texture[49][45] = 0;	doodle_right_transparency_texture[49][46] = 0;	doodle_right_transparency_texture[49][47] = 0;	doodle_right_transparency_texture[49][48] = 0;	doodle_right_transparency_texture[49][49] = 0;	doodle_right_transparency_texture[49][50] = 0;	doodle_right_transparency_texture[49][51] = 0;	doodle_right_transparency_texture[49][52] = 1;	doodle_right_transparency_texture[49][53] = 1;	doodle_right_transparency_texture[49][54] = 1;	doodle_right_transparency_texture[49][55] = 1;	doodle_right_transparency_texture[49][56] = 1;	doodle_right_transparency_texture[49][57] = 1;	doodle_right_transparency_texture[49][58] = 1;	doodle_right_transparency_texture[49][59] = 1;	doodle_right_transparency_texture[49][60] = 1;	doodle_right_transparency_texture[49][61] = 1;	doodle_right_transparency_texture[49][62] = 1;	doodle_right_transparency_texture[49][63] = 1;	doodle_right_transparency_texture[49][64] = 1;	doodle_right_transparency_texture[49][65] = 1;	doodle_right_transparency_texture[49][66] = 1;	doodle_right_transparency_texture[49][67] = 1;	doodle_right_transparency_texture[49][68] = 1;	doodle_right_transparency_texture[49][69] = 1;	doodle_right_transparency_texture[49][70] = 1;	doodle_right_transparency_texture[49][71] = 1;	doodle_right_transparency_texture[49][72] = 1;	doodle_right_transparency_texture[49][73] = 1;	doodle_right_transparency_texture[49][74] = 1;	doodle_right_transparency_texture[49][75] = 1;	doodle_right_transparency_texture[49][76] = 1;	doodle_right_transparency_texture[49][77] = 1;	doodle_right_transparency_texture[49][78] = 1;	doodle_right_transparency_texture[49][79] = 1;	doodle_right_transparency_texture[50][0] = 1;	doodle_right_transparency_texture[50][1] = 1;	doodle_right_transparency_texture[50][2] = 1;	doodle_right_transparency_texture[50][3] = 1;	doodle_right_transparency_texture[50][4] = 0;	doodle_right_transparency_texture[50][5] = 0;	doodle_right_transparency_texture[50][6] = 0;	doodle_right_transparency_texture[50][7] = 0;	doodle_right_transparency_texture[50][8] = 0;	doodle_right_transparency_texture[50][9] = 0;	doodle_right_transparency_texture[50][10] = 0;	doodle_right_transparency_texture[50][11] = 0;	doodle_right_transparency_texture[50][12] = 0;	doodle_right_transparency_texture[50][13] = 0;	doodle_right_transparency_texture[50][14] = 0;	doodle_right_transparency_texture[50][15] = 0;	doodle_right_transparency_texture[50][16] = 0;	doodle_right_transparency_texture[50][17] = 0;	doodle_right_transparency_texture[50][18] = 0;	doodle_right_transparency_texture[50][19] = 0;	doodle_right_transparency_texture[50][20] = 0;	doodle_right_transparency_texture[50][21] = 0;	doodle_right_transparency_texture[50][22] = 0;	doodle_right_transparency_texture[50][23] = 0;	doodle_right_transparency_texture[50][24] = 0;	doodle_right_transparency_texture[50][25] = 0;	doodle_right_transparency_texture[50][26] = 0;	doodle_right_transparency_texture[50][27] = 0;	doodle_right_transparency_texture[50][28] = 0;	doodle_right_transparency_texture[50][29] = 0;	doodle_right_transparency_texture[50][30] = 0;	doodle_right_transparency_texture[50][31] = 0;	doodle_right_transparency_texture[50][32] = 0;	doodle_right_transparency_texture[50][33] = 0;	doodle_right_transparency_texture[50][34] = 0;	doodle_right_transparency_texture[50][35] = 0;	doodle_right_transparency_texture[50][36] = 0;	doodle_right_transparency_texture[50][37] = 0;	doodle_right_transparency_texture[50][38] = 0;	doodle_right_transparency_texture[50][39] = 0;	doodle_right_transparency_texture[50][40] = 0;	doodle_right_transparency_texture[50][41] = 0;	doodle_right_transparency_texture[50][42] = 0;	doodle_right_transparency_texture[50][43] = 0;	doodle_right_transparency_texture[50][44] = 0;	doodle_right_transparency_texture[50][45] = 0;	doodle_right_transparency_texture[50][46] = 0;	doodle_right_transparency_texture[50][47] = 0;	doodle_right_transparency_texture[50][48] = 0;	doodle_right_transparency_texture[50][49] = 0;	doodle_right_transparency_texture[50][50] = 0;	doodle_right_transparency_texture[50][51] = 0;	doodle_right_transparency_texture[50][52] = 1;	doodle_right_transparency_texture[50][53] = 1;	doodle_right_transparency_texture[50][54] = 1;	doodle_right_transparency_texture[50][55] = 1;	doodle_right_transparency_texture[50][56] = 1;	doodle_right_transparency_texture[50][57] = 1;	doodle_right_transparency_texture[50][58] = 1;	doodle_right_transparency_texture[50][59] = 1;	doodle_right_transparency_texture[50][60] = 1;	doodle_right_transparency_texture[50][61] = 1;	doodle_right_transparency_texture[50][62] = 1;	doodle_right_transparency_texture[50][63] = 1;	doodle_right_transparency_texture[50][64] = 1;	doodle_right_transparency_texture[50][65] = 1;	doodle_right_transparency_texture[50][66] = 1;	doodle_right_transparency_texture[50][67] = 1;	doodle_right_transparency_texture[50][68] = 1;	doodle_right_transparency_texture[50][69] = 1;	doodle_right_transparency_texture[50][70] = 1;	doodle_right_transparency_texture[50][71] = 1;	doodle_right_transparency_texture[50][72] = 1;	doodle_right_transparency_texture[50][73] = 1;	doodle_right_transparency_texture[50][74] = 1;	doodle_right_transparency_texture[50][75] = 1;	doodle_right_transparency_texture[50][76] = 1;	doodle_right_transparency_texture[50][77] = 1;	doodle_right_transparency_texture[50][78] = 1;	doodle_right_transparency_texture[50][79] = 1;	doodle_right_transparency_texture[51][0] = 1;	doodle_right_transparency_texture[51][1] = 1;	doodle_right_transparency_texture[51][2] = 1;	doodle_right_transparency_texture[51][3] = 1;	doodle_right_transparency_texture[51][4] = 0;	doodle_right_transparency_texture[51][5] = 0;	doodle_right_transparency_texture[51][6] = 0;	doodle_right_transparency_texture[51][7] = 0;	doodle_right_transparency_texture[51][8] = 0;	doodle_right_transparency_texture[51][9] = 0;	doodle_right_transparency_texture[51][10] = 0;	doodle_right_transparency_texture[51][11] = 0;	doodle_right_transparency_texture[51][12] = 0;	doodle_right_transparency_texture[51][13] = 0;	doodle_right_transparency_texture[51][14] = 0;	doodle_right_transparency_texture[51][15] = 0;	doodle_right_transparency_texture[51][16] = 0;	doodle_right_transparency_texture[51][17] = 0;	doodle_right_transparency_texture[51][18] = 0;	doodle_right_transparency_texture[51][19] = 0;	doodle_right_transparency_texture[51][20] = 0;	doodle_right_transparency_texture[51][21] = 0;	doodle_right_transparency_texture[51][22] = 0;	doodle_right_transparency_texture[51][23] = 0;	doodle_right_transparency_texture[51][24] = 0;	doodle_right_transparency_texture[51][25] = 0;	doodle_right_transparency_texture[51][26] = 0;	doodle_right_transparency_texture[51][27] = 0;	doodle_right_transparency_texture[51][28] = 0;	doodle_right_transparency_texture[51][29] = 0;	doodle_right_transparency_texture[51][30] = 0;	doodle_right_transparency_texture[51][31] = 0;	doodle_right_transparency_texture[51][32] = 0;	doodle_right_transparency_texture[51][33] = 0;	doodle_right_transparency_texture[51][34] = 0;	doodle_right_transparency_texture[51][35] = 0;	doodle_right_transparency_texture[51][36] = 0;	doodle_right_transparency_texture[51][37] = 0;	doodle_right_transparency_texture[51][38] = 0;	doodle_right_transparency_texture[51][39] = 0;	doodle_right_transparency_texture[51][40] = 0;	doodle_right_transparency_texture[51][41] = 0;	doodle_right_transparency_texture[51][42] = 0;	doodle_right_transparency_texture[51][43] = 0;	doodle_right_transparency_texture[51][44] = 0;	doodle_right_transparency_texture[51][45] = 0;	doodle_right_transparency_texture[51][46] = 0;	doodle_right_transparency_texture[51][47] = 0;	doodle_right_transparency_texture[51][48] = 0;	doodle_right_transparency_texture[51][49] = 0;	doodle_right_transparency_texture[51][50] = 0;	doodle_right_transparency_texture[51][51] = 0;	doodle_right_transparency_texture[51][52] = 1;	doodle_right_transparency_texture[51][53] = 1;	doodle_right_transparency_texture[51][54] = 1;	doodle_right_transparency_texture[51][55] = 1;	doodle_right_transparency_texture[51][56] = 1;	doodle_right_transparency_texture[51][57] = 1;	doodle_right_transparency_texture[51][58] = 1;	doodle_right_transparency_texture[51][59] = 1;	doodle_right_transparency_texture[51][60] = 1;	doodle_right_transparency_texture[51][61] = 1;	doodle_right_transparency_texture[51][62] = 1;	doodle_right_transparency_texture[51][63] = 1;	doodle_right_transparency_texture[51][64] = 1;	doodle_right_transparency_texture[51][65] = 1;	doodle_right_transparency_texture[51][66] = 1;	doodle_right_transparency_texture[51][67] = 1;	doodle_right_transparency_texture[51][68] = 1;	doodle_right_transparency_texture[51][69] = 1;	doodle_right_transparency_texture[51][70] = 1;	doodle_right_transparency_texture[51][71] = 1;	doodle_right_transparency_texture[51][72] = 1;	doodle_right_transparency_texture[51][73] = 1;	doodle_right_transparency_texture[51][74] = 1;	doodle_right_transparency_texture[51][75] = 1;	doodle_right_transparency_texture[51][76] = 1;	doodle_right_transparency_texture[51][77] = 1;	doodle_right_transparency_texture[51][78] = 1;	doodle_right_transparency_texture[51][79] = 1;	doodle_right_transparency_texture[52][0] = 1;	doodle_right_transparency_texture[52][1] = 1;	doodle_right_transparency_texture[52][2] = 1;	doodle_right_transparency_texture[52][3] = 1;	doodle_right_transparency_texture[52][4] = 0;	doodle_right_transparency_texture[52][5] = 0;	doodle_right_transparency_texture[52][6] = 0;	doodle_right_transparency_texture[52][7] = 0;	doodle_right_transparency_texture[52][8] = 0;	doodle_right_transparency_texture[52][9] = 0;	doodle_right_transparency_texture[52][10] = 0;	doodle_right_transparency_texture[52][11] = 0;	doodle_right_transparency_texture[52][12] = 0;	doodle_right_transparency_texture[52][13] = 0;	doodle_right_transparency_texture[52][14] = 0;	doodle_right_transparency_texture[52][15] = 0;	doodle_right_transparency_texture[52][16] = 0;	doodle_right_transparency_texture[52][17] = 0;	doodle_right_transparency_texture[52][18] = 0;	doodle_right_transparency_texture[52][19] = 0;	doodle_right_transparency_texture[52][20] = 0;	doodle_right_transparency_texture[52][21] = 0;	doodle_right_transparency_texture[52][22] = 0;	doodle_right_transparency_texture[52][23] = 0;	doodle_right_transparency_texture[52][24] = 0;	doodle_right_transparency_texture[52][25] = 0;	doodle_right_transparency_texture[52][26] = 0;	doodle_right_transparency_texture[52][27] = 0;	doodle_right_transparency_texture[52][28] = 0;	doodle_right_transparency_texture[52][29] = 0;	doodle_right_transparency_texture[52][30] = 0;	doodle_right_transparency_texture[52][31] = 0;	doodle_right_transparency_texture[52][32] = 0;	doodle_right_transparency_texture[52][33] = 0;	doodle_right_transparency_texture[52][34] = 0;	doodle_right_transparency_texture[52][35] = 0;	doodle_right_transparency_texture[52][36] = 0;	doodle_right_transparency_texture[52][37] = 0;	doodle_right_transparency_texture[52][38] = 0;	doodle_right_transparency_texture[52][39] = 0;	doodle_right_transparency_texture[52][40] = 0;	doodle_right_transparency_texture[52][41] = 0;	doodle_right_transparency_texture[52][42] = 0;	doodle_right_transparency_texture[52][43] = 0;	doodle_right_transparency_texture[52][44] = 0;	doodle_right_transparency_texture[52][45] = 0;	doodle_right_transparency_texture[52][46] = 0;	doodle_right_transparency_texture[52][47] = 0;	doodle_right_transparency_texture[52][48] = 0;	doodle_right_transparency_texture[52][49] = 0;	doodle_right_transparency_texture[52][50] = 0;	doodle_right_transparency_texture[52][51] = 0;	doodle_right_transparency_texture[52][52] = 1;	doodle_right_transparency_texture[52][53] = 1;	doodle_right_transparency_texture[52][54] = 1;	doodle_right_transparency_texture[52][55] = 1;	doodle_right_transparency_texture[52][56] = 1;	doodle_right_transparency_texture[52][57] = 1;	doodle_right_transparency_texture[52][58] = 1;	doodle_right_transparency_texture[52][59] = 1;	doodle_right_transparency_texture[52][60] = 1;	doodle_right_transparency_texture[52][61] = 1;	doodle_right_transparency_texture[52][62] = 1;	doodle_right_transparency_texture[52][63] = 1;	doodle_right_transparency_texture[52][64] = 1;	doodle_right_transparency_texture[52][65] = 1;	doodle_right_transparency_texture[52][66] = 1;	doodle_right_transparency_texture[52][67] = 1;	doodle_right_transparency_texture[52][68] = 1;	doodle_right_transparency_texture[52][69] = 1;	doodle_right_transparency_texture[52][70] = 1;	doodle_right_transparency_texture[52][71] = 1;	doodle_right_transparency_texture[52][72] = 1;	doodle_right_transparency_texture[52][73] = 1;	doodle_right_transparency_texture[52][74] = 1;	doodle_right_transparency_texture[52][75] = 1;	doodle_right_transparency_texture[52][76] = 1;	doodle_right_transparency_texture[52][77] = 1;	doodle_right_transparency_texture[52][78] = 1;	doodle_right_transparency_texture[52][79] = 1;	doodle_right_transparency_texture[53][0] = 1;	doodle_right_transparency_texture[53][1] = 1;	doodle_right_transparency_texture[53][2] = 1;	doodle_right_transparency_texture[53][3] = 1;	doodle_right_transparency_texture[53][4] = 0;	doodle_right_transparency_texture[53][5] = 0;	doodle_right_transparency_texture[53][6] = 0;	doodle_right_transparency_texture[53][7] = 0;	doodle_right_transparency_texture[53][8] = 0;	doodle_right_transparency_texture[53][9] = 0;	doodle_right_transparency_texture[53][10] = 0;	doodle_right_transparency_texture[53][11] = 0;	doodle_right_transparency_texture[53][12] = 0;	doodle_right_transparency_texture[53][13] = 0;	doodle_right_transparency_texture[53][14] = 0;	doodle_right_transparency_texture[53][15] = 0;	doodle_right_transparency_texture[53][16] = 0;	doodle_right_transparency_texture[53][17] = 0;	doodle_right_transparency_texture[53][18] = 0;	doodle_right_transparency_texture[53][19] = 0;	doodle_right_transparency_texture[53][20] = 0;	doodle_right_transparency_texture[53][21] = 0;	doodle_right_transparency_texture[53][22] = 0;	doodle_right_transparency_texture[53][23] = 0;	doodle_right_transparency_texture[53][24] = 0;	doodle_right_transparency_texture[53][25] = 0;	doodle_right_transparency_texture[53][26] = 0;	doodle_right_transparency_texture[53][27] = 0;	doodle_right_transparency_texture[53][28] = 0;	doodle_right_transparency_texture[53][29] = 0;	doodle_right_transparency_texture[53][30] = 0;	doodle_right_transparency_texture[53][31] = 0;	doodle_right_transparency_texture[53][32] = 0;	doodle_right_transparency_texture[53][33] = 0;	doodle_right_transparency_texture[53][34] = 0;	doodle_right_transparency_texture[53][35] = 0;	doodle_right_transparency_texture[53][36] = 0;	doodle_right_transparency_texture[53][37] = 0;	doodle_right_transparency_texture[53][38] = 0;	doodle_right_transparency_texture[53][39] = 0;	doodle_right_transparency_texture[53][40] = 0;	doodle_right_transparency_texture[53][41] = 0;	doodle_right_transparency_texture[53][42] = 0;	doodle_right_transparency_texture[53][43] = 0;	doodle_right_transparency_texture[53][44] = 0;	doodle_right_transparency_texture[53][45] = 0;	doodle_right_transparency_texture[53][46] = 0;	doodle_right_transparency_texture[53][47] = 0;	doodle_right_transparency_texture[53][48] = 0;	doodle_right_transparency_texture[53][49] = 0;	doodle_right_transparency_texture[53][50] = 0;	doodle_right_transparency_texture[53][51] = 0;	doodle_right_transparency_texture[53][52] = 1;	doodle_right_transparency_texture[53][53] = 1;	doodle_right_transparency_texture[53][54] = 1;	doodle_right_transparency_texture[53][55] = 1;	doodle_right_transparency_texture[53][56] = 1;	doodle_right_transparency_texture[53][57] = 1;	doodle_right_transparency_texture[53][58] = 1;	doodle_right_transparency_texture[53][59] = 1;	doodle_right_transparency_texture[53][60] = 1;	doodle_right_transparency_texture[53][61] = 1;	doodle_right_transparency_texture[53][62] = 1;	doodle_right_transparency_texture[53][63] = 1;	doodle_right_transparency_texture[53][64] = 1;	doodle_right_transparency_texture[53][65] = 1;	doodle_right_transparency_texture[53][66] = 1;	doodle_right_transparency_texture[53][67] = 1;	doodle_right_transparency_texture[53][68] = 1;	doodle_right_transparency_texture[53][69] = 1;	doodle_right_transparency_texture[53][70] = 1;	doodle_right_transparency_texture[53][71] = 1;	doodle_right_transparency_texture[53][72] = 1;	doodle_right_transparency_texture[53][73] = 1;	doodle_right_transparency_texture[53][74] = 1;	doodle_right_transparency_texture[53][75] = 1;	doodle_right_transparency_texture[53][76] = 1;	doodle_right_transparency_texture[53][77] = 1;	doodle_right_transparency_texture[53][78] = 1;	doodle_right_transparency_texture[53][79] = 1;	doodle_right_transparency_texture[54][0] = 1;	doodle_right_transparency_texture[54][1] = 1;	doodle_right_transparency_texture[54][2] = 1;	doodle_right_transparency_texture[54][3] = 1;	doodle_right_transparency_texture[54][4] = 0;	doodle_right_transparency_texture[54][5] = 0;	doodle_right_transparency_texture[54][6] = 0;	doodle_right_transparency_texture[54][7] = 0;	doodle_right_transparency_texture[54][8] = 0;	doodle_right_transparency_texture[54][9] = 0;	doodle_right_transparency_texture[54][10] = 0;	doodle_right_transparency_texture[54][11] = 0;	doodle_right_transparency_texture[54][12] = 0;	doodle_right_transparency_texture[54][13] = 0;	doodle_right_transparency_texture[54][14] = 0;	doodle_right_transparency_texture[54][15] = 0;	doodle_right_transparency_texture[54][16] = 0;	doodle_right_transparency_texture[54][17] = 0;	doodle_right_transparency_texture[54][18] = 0;	doodle_right_transparency_texture[54][19] = 0;	doodle_right_transparency_texture[54][20] = 0;	doodle_right_transparency_texture[54][21] = 0;	doodle_right_transparency_texture[54][22] = 0;	doodle_right_transparency_texture[54][23] = 0;	doodle_right_transparency_texture[54][24] = 0;	doodle_right_transparency_texture[54][25] = 0;	doodle_right_transparency_texture[54][26] = 0;	doodle_right_transparency_texture[54][27] = 0;	doodle_right_transparency_texture[54][28] = 0;	doodle_right_transparency_texture[54][29] = 0;	doodle_right_transparency_texture[54][30] = 0;	doodle_right_transparency_texture[54][31] = 0;	doodle_right_transparency_texture[54][32] = 0;	doodle_right_transparency_texture[54][33] = 0;	doodle_right_transparency_texture[54][34] = 0;	doodle_right_transparency_texture[54][35] = 0;	doodle_right_transparency_texture[54][36] = 0;	doodle_right_transparency_texture[54][37] = 0;	doodle_right_transparency_texture[54][38] = 0;	doodle_right_transparency_texture[54][39] = 0;	doodle_right_transparency_texture[54][40] = 0;	doodle_right_transparency_texture[54][41] = 0;	doodle_right_transparency_texture[54][42] = 0;	doodle_right_transparency_texture[54][43] = 0;	doodle_right_transparency_texture[54][44] = 0;	doodle_right_transparency_texture[54][45] = 0;	doodle_right_transparency_texture[54][46] = 0;	doodle_right_transparency_texture[54][47] = 0;	doodle_right_transparency_texture[54][48] = 0;	doodle_right_transparency_texture[54][49] = 0;	doodle_right_transparency_texture[54][50] = 0;	doodle_right_transparency_texture[54][51] = 0;	doodle_right_transparency_texture[54][52] = 1;	doodle_right_transparency_texture[54][53] = 1;	doodle_right_transparency_texture[54][54] = 1;	doodle_right_transparency_texture[54][55] = 1;	doodle_right_transparency_texture[54][56] = 1;	doodle_right_transparency_texture[54][57] = 1;	doodle_right_transparency_texture[54][58] = 1;	doodle_right_transparency_texture[54][59] = 1;	doodle_right_transparency_texture[54][60] = 1;	doodle_right_transparency_texture[54][61] = 1;	doodle_right_transparency_texture[54][62] = 1;	doodle_right_transparency_texture[54][63] = 1;	doodle_right_transparency_texture[54][64] = 1;	doodle_right_transparency_texture[54][65] = 1;	doodle_right_transparency_texture[54][66] = 1;	doodle_right_transparency_texture[54][67] = 1;	doodle_right_transparency_texture[54][68] = 1;	doodle_right_transparency_texture[54][69] = 1;	doodle_right_transparency_texture[54][70] = 1;	doodle_right_transparency_texture[54][71] = 1;	doodle_right_transparency_texture[54][72] = 1;	doodle_right_transparency_texture[54][73] = 1;	doodle_right_transparency_texture[54][74] = 1;	doodle_right_transparency_texture[54][75] = 1;	doodle_right_transparency_texture[54][76] = 1;	doodle_right_transparency_texture[54][77] = 1;	doodle_right_transparency_texture[54][78] = 1;	doodle_right_transparency_texture[54][79] = 1;	doodle_right_transparency_texture[55][0] = 1;	doodle_right_transparency_texture[55][1] = 1;	doodle_right_transparency_texture[55][2] = 1;	doodle_right_transparency_texture[55][3] = 1;	doodle_right_transparency_texture[55][4] = 0;	doodle_right_transparency_texture[55][5] = 0;	doodle_right_transparency_texture[55][6] = 0;	doodle_right_transparency_texture[55][7] = 0;	doodle_right_transparency_texture[55][8] = 0;	doodle_right_transparency_texture[55][9] = 0;	doodle_right_transparency_texture[55][10] = 0;	doodle_right_transparency_texture[55][11] = 0;	doodle_right_transparency_texture[55][12] = 0;	doodle_right_transparency_texture[55][13] = 0;	doodle_right_transparency_texture[55][14] = 0;	doodle_right_transparency_texture[55][15] = 0;	doodle_right_transparency_texture[55][16] = 0;	doodle_right_transparency_texture[55][17] = 0;	doodle_right_transparency_texture[55][18] = 0;	doodle_right_transparency_texture[55][19] = 0;	doodle_right_transparency_texture[55][20] = 0;	doodle_right_transparency_texture[55][21] = 0;	doodle_right_transparency_texture[55][22] = 0;	doodle_right_transparency_texture[55][23] = 0;	doodle_right_transparency_texture[55][24] = 0;	doodle_right_transparency_texture[55][25] = 0;	doodle_right_transparency_texture[55][26] = 0;	doodle_right_transparency_texture[55][27] = 0;	doodle_right_transparency_texture[55][28] = 0;	doodle_right_transparency_texture[55][29] = 0;	doodle_right_transparency_texture[55][30] = 0;	doodle_right_transparency_texture[55][31] = 0;	doodle_right_transparency_texture[55][32] = 0;	doodle_right_transparency_texture[55][33] = 0;	doodle_right_transparency_texture[55][34] = 0;	doodle_right_transparency_texture[55][35] = 0;	doodle_right_transparency_texture[55][36] = 0;	doodle_right_transparency_texture[55][37] = 0;	doodle_right_transparency_texture[55][38] = 0;	doodle_right_transparency_texture[55][39] = 0;	doodle_right_transparency_texture[55][40] = 0;	doodle_right_transparency_texture[55][41] = 0;	doodle_right_transparency_texture[55][42] = 0;	doodle_right_transparency_texture[55][43] = 0;	doodle_right_transparency_texture[55][44] = 0;	doodle_right_transparency_texture[55][45] = 0;	doodle_right_transparency_texture[55][46] = 0;	doodle_right_transparency_texture[55][47] = 0;	doodle_right_transparency_texture[55][48] = 0;	doodle_right_transparency_texture[55][49] = 0;	doodle_right_transparency_texture[55][50] = 0;	doodle_right_transparency_texture[55][51] = 0;	doodle_right_transparency_texture[55][52] = 1;	doodle_right_transparency_texture[55][53] = 1;	doodle_right_transparency_texture[55][54] = 1;	doodle_right_transparency_texture[55][55] = 1;	doodle_right_transparency_texture[55][56] = 1;	doodle_right_transparency_texture[55][57] = 1;	doodle_right_transparency_texture[55][58] = 1;	doodle_right_transparency_texture[55][59] = 1;	doodle_right_transparency_texture[55][60] = 1;	doodle_right_transparency_texture[55][61] = 1;	doodle_right_transparency_texture[55][62] = 1;	doodle_right_transparency_texture[55][63] = 1;	doodle_right_transparency_texture[55][64] = 1;	doodle_right_transparency_texture[55][65] = 1;	doodle_right_transparency_texture[55][66] = 1;	doodle_right_transparency_texture[55][67] = 1;	doodle_right_transparency_texture[55][68] = 1;	doodle_right_transparency_texture[55][69] = 1;	doodle_right_transparency_texture[55][70] = 1;	doodle_right_transparency_texture[55][71] = 1;	doodle_right_transparency_texture[55][72] = 1;	doodle_right_transparency_texture[55][73] = 1;	doodle_right_transparency_texture[55][74] = 1;	doodle_right_transparency_texture[55][75] = 1;	doodle_right_transparency_texture[55][76] = 1;	doodle_right_transparency_texture[55][77] = 1;	doodle_right_transparency_texture[55][78] = 1;	doodle_right_transparency_texture[55][79] = 1;	doodle_right_transparency_texture[56][0] = 1;	doodle_right_transparency_texture[56][1] = 1;	doodle_right_transparency_texture[56][2] = 1;	doodle_right_transparency_texture[56][3] = 1;	doodle_right_transparency_texture[56][4] = 0;	doodle_right_transparency_texture[56][5] = 0;	doodle_right_transparency_texture[56][6] = 0;	doodle_right_transparency_texture[56][7] = 0;	doodle_right_transparency_texture[56][8] = 0;	doodle_right_transparency_texture[56][9] = 0;	doodle_right_transparency_texture[56][10] = 0;	doodle_right_transparency_texture[56][11] = 0;	doodle_right_transparency_texture[56][12] = 0;	doodle_right_transparency_texture[56][13] = 0;	doodle_right_transparency_texture[56][14] = 0;	doodle_right_transparency_texture[56][15] = 0;	doodle_right_transparency_texture[56][16] = 0;	doodle_right_transparency_texture[56][17] = 0;	doodle_right_transparency_texture[56][18] = 0;	doodle_right_transparency_texture[56][19] = 0;	doodle_right_transparency_texture[56][20] = 0;	doodle_right_transparency_texture[56][21] = 0;	doodle_right_transparency_texture[56][22] = 0;	doodle_right_transparency_texture[56][23] = 0;	doodle_right_transparency_texture[56][24] = 0;	doodle_right_transparency_texture[56][25] = 0;	doodle_right_transparency_texture[56][26] = 0;	doodle_right_transparency_texture[56][27] = 0;	doodle_right_transparency_texture[56][28] = 0;	doodle_right_transparency_texture[56][29] = 0;	doodle_right_transparency_texture[56][30] = 0;	doodle_right_transparency_texture[56][31] = 0;	doodle_right_transparency_texture[56][32] = 0;	doodle_right_transparency_texture[56][33] = 0;	doodle_right_transparency_texture[56][34] = 0;	doodle_right_transparency_texture[56][35] = 0;	doodle_right_transparency_texture[56][36] = 0;	doodle_right_transparency_texture[56][37] = 0;	doodle_right_transparency_texture[56][38] = 0;	doodle_right_transparency_texture[56][39] = 0;	doodle_right_transparency_texture[56][40] = 0;	doodle_right_transparency_texture[56][41] = 0;	doodle_right_transparency_texture[56][42] = 0;	doodle_right_transparency_texture[56][43] = 0;	doodle_right_transparency_texture[56][44] = 0;	doodle_right_transparency_texture[56][45] = 0;	doodle_right_transparency_texture[56][46] = 0;	doodle_right_transparency_texture[56][47] = 0;	doodle_right_transparency_texture[56][48] = 0;	doodle_right_transparency_texture[56][49] = 0;	doodle_right_transparency_texture[56][50] = 0;	doodle_right_transparency_texture[56][51] = 0;	doodle_right_transparency_texture[56][52] = 1;	doodle_right_transparency_texture[56][53] = 1;	doodle_right_transparency_texture[56][54] = 1;	doodle_right_transparency_texture[56][55] = 1;	doodle_right_transparency_texture[56][56] = 1;	doodle_right_transparency_texture[56][57] = 1;	doodle_right_transparency_texture[56][58] = 1;	doodle_right_transparency_texture[56][59] = 1;	doodle_right_transparency_texture[56][60] = 1;	doodle_right_transparency_texture[56][61] = 1;	doodle_right_transparency_texture[56][62] = 1;	doodle_right_transparency_texture[56][63] = 1;	doodle_right_transparency_texture[56][64] = 1;	doodle_right_transparency_texture[56][65] = 1;	doodle_right_transparency_texture[56][66] = 1;	doodle_right_transparency_texture[56][67] = 1;	doodle_right_transparency_texture[56][68] = 1;	doodle_right_transparency_texture[56][69] = 1;	doodle_right_transparency_texture[56][70] = 1;	doodle_right_transparency_texture[56][71] = 1;	doodle_right_transparency_texture[56][72] = 1;	doodle_right_transparency_texture[56][73] = 1;	doodle_right_transparency_texture[56][74] = 1;	doodle_right_transparency_texture[56][75] = 1;	doodle_right_transparency_texture[56][76] = 1;	doodle_right_transparency_texture[56][77] = 1;	doodle_right_transparency_texture[56][78] = 1;	doodle_right_transparency_texture[56][79] = 1;	doodle_right_transparency_texture[57][0] = 1;	doodle_right_transparency_texture[57][1] = 1;	doodle_right_transparency_texture[57][2] = 1;	doodle_right_transparency_texture[57][3] = 1;	doodle_right_transparency_texture[57][4] = 0;	doodle_right_transparency_texture[57][5] = 0;	doodle_right_transparency_texture[57][6] = 0;	doodle_right_transparency_texture[57][7] = 0;	doodle_right_transparency_texture[57][8] = 0;	doodle_right_transparency_texture[57][9] = 0;	doodle_right_transparency_texture[57][10] = 0;	doodle_right_transparency_texture[57][11] = 0;	doodle_right_transparency_texture[57][12] = 0;	doodle_right_transparency_texture[57][13] = 0;	doodle_right_transparency_texture[57][14] = 0;	doodle_right_transparency_texture[57][15] = 0;	doodle_right_transparency_texture[57][16] = 0;	doodle_right_transparency_texture[57][17] = 0;	doodle_right_transparency_texture[57][18] = 0;	doodle_right_transparency_texture[57][19] = 0;	doodle_right_transparency_texture[57][20] = 0;	doodle_right_transparency_texture[57][21] = 0;	doodle_right_transparency_texture[57][22] = 0;	doodle_right_transparency_texture[57][23] = 0;	doodle_right_transparency_texture[57][24] = 0;	doodle_right_transparency_texture[57][25] = 0;	doodle_right_transparency_texture[57][26] = 0;	doodle_right_transparency_texture[57][27] = 0;	doodle_right_transparency_texture[57][28] = 0;	doodle_right_transparency_texture[57][29] = 0;	doodle_right_transparency_texture[57][30] = 0;	doodle_right_transparency_texture[57][31] = 0;	doodle_right_transparency_texture[57][32] = 0;	doodle_right_transparency_texture[57][33] = 0;	doodle_right_transparency_texture[57][34] = 0;	doodle_right_transparency_texture[57][35] = 0;	doodle_right_transparency_texture[57][36] = 0;	doodle_right_transparency_texture[57][37] = 0;	doodle_right_transparency_texture[57][38] = 0;	doodle_right_transparency_texture[57][39] = 0;	doodle_right_transparency_texture[57][40] = 0;	doodle_right_transparency_texture[57][41] = 0;	doodle_right_transparency_texture[57][42] = 0;	doodle_right_transparency_texture[57][43] = 0;	doodle_right_transparency_texture[57][44] = 0;	doodle_right_transparency_texture[57][45] = 0;	doodle_right_transparency_texture[57][46] = 0;	doodle_right_transparency_texture[57][47] = 0;	doodle_right_transparency_texture[57][48] = 0;	doodle_right_transparency_texture[57][49] = 0;	doodle_right_transparency_texture[57][50] = 0;	doodle_right_transparency_texture[57][51] = 0;	doodle_right_transparency_texture[57][52] = 1;	doodle_right_transparency_texture[57][53] = 1;	doodle_right_transparency_texture[57][54] = 1;	doodle_right_transparency_texture[57][55] = 1;	doodle_right_transparency_texture[57][56] = 1;	doodle_right_transparency_texture[57][57] = 1;	doodle_right_transparency_texture[57][58] = 1;	doodle_right_transparency_texture[57][59] = 1;	doodle_right_transparency_texture[57][60] = 1;	doodle_right_transparency_texture[57][61] = 1;	doodle_right_transparency_texture[57][62] = 1;	doodle_right_transparency_texture[57][63] = 1;	doodle_right_transparency_texture[57][64] = 1;	doodle_right_transparency_texture[57][65] = 1;	doodle_right_transparency_texture[57][66] = 1;	doodle_right_transparency_texture[57][67] = 1;	doodle_right_transparency_texture[57][68] = 1;	doodle_right_transparency_texture[57][69] = 1;	doodle_right_transparency_texture[57][70] = 1;	doodle_right_transparency_texture[57][71] = 1;	doodle_right_transparency_texture[57][72] = 1;	doodle_right_transparency_texture[57][73] = 1;	doodle_right_transparency_texture[57][74] = 1;	doodle_right_transparency_texture[57][75] = 1;	doodle_right_transparency_texture[57][76] = 1;	doodle_right_transparency_texture[57][77] = 1;	doodle_right_transparency_texture[57][78] = 1;	doodle_right_transparency_texture[57][79] = 1;	doodle_right_transparency_texture[58][0] = 1;	doodle_right_transparency_texture[58][1] = 1;	doodle_right_transparency_texture[58][2] = 1;	doodle_right_transparency_texture[58][3] = 1;	doodle_right_transparency_texture[58][4] = 0;	doodle_right_transparency_texture[58][5] = 0;	doodle_right_transparency_texture[58][6] = 0;	doodle_right_transparency_texture[58][7] = 0;	doodle_right_transparency_texture[58][8] = 0;	doodle_right_transparency_texture[58][9] = 0;	doodle_right_transparency_texture[58][10] = 0;	doodle_right_transparency_texture[58][11] = 0;	doodle_right_transparency_texture[58][12] = 0;	doodle_right_transparency_texture[58][13] = 0;	doodle_right_transparency_texture[58][14] = 0;	doodle_right_transparency_texture[58][15] = 0;	doodle_right_transparency_texture[58][16] = 0;	doodle_right_transparency_texture[58][17] = 0;	doodle_right_transparency_texture[58][18] = 0;	doodle_right_transparency_texture[58][19] = 0;	doodle_right_transparency_texture[58][20] = 0;	doodle_right_transparency_texture[58][21] = 0;	doodle_right_transparency_texture[58][22] = 0;	doodle_right_transparency_texture[58][23] = 0;	doodle_right_transparency_texture[58][24] = 0;	doodle_right_transparency_texture[58][25] = 0;	doodle_right_transparency_texture[58][26] = 0;	doodle_right_transparency_texture[58][27] = 0;	doodle_right_transparency_texture[58][28] = 0;	doodle_right_transparency_texture[58][29] = 0;	doodle_right_transparency_texture[58][30] = 0;	doodle_right_transparency_texture[58][31] = 0;	doodle_right_transparency_texture[58][32] = 0;	doodle_right_transparency_texture[58][33] = 0;	doodle_right_transparency_texture[58][34] = 0;	doodle_right_transparency_texture[58][35] = 0;	doodle_right_transparency_texture[58][36] = 0;	doodle_right_transparency_texture[58][37] = 0;	doodle_right_transparency_texture[58][38] = 0;	doodle_right_transparency_texture[58][39] = 0;	doodle_right_transparency_texture[58][40] = 0;	doodle_right_transparency_texture[58][41] = 0;	doodle_right_transparency_texture[58][42] = 0;	doodle_right_transparency_texture[58][43] = 0;	doodle_right_transparency_texture[58][44] = 0;	doodle_right_transparency_texture[58][45] = 0;	doodle_right_transparency_texture[58][46] = 0;	doodle_right_transparency_texture[58][47] = 0;	doodle_right_transparency_texture[58][48] = 0;	doodle_right_transparency_texture[58][49] = 0;	doodle_right_transparency_texture[58][50] = 0;	doodle_right_transparency_texture[58][51] = 0;	doodle_right_transparency_texture[58][52] = 1;	doodle_right_transparency_texture[58][53] = 1;	doodle_right_transparency_texture[58][54] = 1;	doodle_right_transparency_texture[58][55] = 1;	doodle_right_transparency_texture[58][56] = 1;	doodle_right_transparency_texture[58][57] = 1;	doodle_right_transparency_texture[58][58] = 1;	doodle_right_transparency_texture[58][59] = 1;	doodle_right_transparency_texture[58][60] = 1;	doodle_right_transparency_texture[58][61] = 1;	doodle_right_transparency_texture[58][62] = 1;	doodle_right_transparency_texture[58][63] = 1;	doodle_right_transparency_texture[58][64] = 1;	doodle_right_transparency_texture[58][65] = 1;	doodle_right_transparency_texture[58][66] = 1;	doodle_right_transparency_texture[58][67] = 1;	doodle_right_transparency_texture[58][68] = 1;	doodle_right_transparency_texture[58][69] = 1;	doodle_right_transparency_texture[58][70] = 1;	doodle_right_transparency_texture[58][71] = 1;	doodle_right_transparency_texture[58][72] = 1;	doodle_right_transparency_texture[58][73] = 1;	doodle_right_transparency_texture[58][74] = 1;	doodle_right_transparency_texture[58][75] = 1;	doodle_right_transparency_texture[58][76] = 1;	doodle_right_transparency_texture[58][77] = 1;	doodle_right_transparency_texture[58][78] = 1;	doodle_right_transparency_texture[58][79] = 1;	doodle_right_transparency_texture[59][0] = 1;	doodle_right_transparency_texture[59][1] = 1;	doodle_right_transparency_texture[59][2] = 1;	doodle_right_transparency_texture[59][3] = 1;	doodle_right_transparency_texture[59][4] = 0;	doodle_right_transparency_texture[59][5] = 0;	doodle_right_transparency_texture[59][6] = 0;	doodle_right_transparency_texture[59][7] = 0;	doodle_right_transparency_texture[59][8] = 0;	doodle_right_transparency_texture[59][9] = 0;	doodle_right_transparency_texture[59][10] = 0;	doodle_right_transparency_texture[59][11] = 0;	doodle_right_transparency_texture[59][12] = 0;	doodle_right_transparency_texture[59][13] = 0;	doodle_right_transparency_texture[59][14] = 0;	doodle_right_transparency_texture[59][15] = 0;	doodle_right_transparency_texture[59][16] = 0;	doodle_right_transparency_texture[59][17] = 0;	doodle_right_transparency_texture[59][18] = 0;	doodle_right_transparency_texture[59][19] = 0;	doodle_right_transparency_texture[59][20] = 0;	doodle_right_transparency_texture[59][21] = 0;	doodle_right_transparency_texture[59][22] = 0;	doodle_right_transparency_texture[59][23] = 0;	doodle_right_transparency_texture[59][24] = 0;	doodle_right_transparency_texture[59][25] = 0;	doodle_right_transparency_texture[59][26] = 0;	doodle_right_transparency_texture[59][27] = 0;	doodle_right_transparency_texture[59][28] = 0;	doodle_right_transparency_texture[59][29] = 0;	doodle_right_transparency_texture[59][30] = 0;	doodle_right_transparency_texture[59][31] = 0;	doodle_right_transparency_texture[59][32] = 0;	doodle_right_transparency_texture[59][33] = 0;	doodle_right_transparency_texture[59][34] = 0;	doodle_right_transparency_texture[59][35] = 0;	doodle_right_transparency_texture[59][36] = 0;	doodle_right_transparency_texture[59][37] = 0;	doodle_right_transparency_texture[59][38] = 0;	doodle_right_transparency_texture[59][39] = 0;	doodle_right_transparency_texture[59][40] = 0;	doodle_right_transparency_texture[59][41] = 0;	doodle_right_transparency_texture[59][42] = 0;	doodle_right_transparency_texture[59][43] = 0;	doodle_right_transparency_texture[59][44] = 0;	doodle_right_transparency_texture[59][45] = 0;	doodle_right_transparency_texture[59][46] = 0;	doodle_right_transparency_texture[59][47] = 0;	doodle_right_transparency_texture[59][48] = 0;	doodle_right_transparency_texture[59][49] = 0;	doodle_right_transparency_texture[59][50] = 0;	doodle_right_transparency_texture[59][51] = 0;	doodle_right_transparency_texture[59][52] = 1;	doodle_right_transparency_texture[59][53] = 1;	doodle_right_transparency_texture[59][54] = 1;	doodle_right_transparency_texture[59][55] = 1;	doodle_right_transparency_texture[59][56] = 1;	doodle_right_transparency_texture[59][57] = 1;	doodle_right_transparency_texture[59][58] = 1;	doodle_right_transparency_texture[59][59] = 1;	doodle_right_transparency_texture[59][60] = 1;	doodle_right_transparency_texture[59][61] = 1;	doodle_right_transparency_texture[59][62] = 1;	doodle_right_transparency_texture[59][63] = 1;	doodle_right_transparency_texture[59][64] = 1;	doodle_right_transparency_texture[59][65] = 1;	doodle_right_transparency_texture[59][66] = 1;	doodle_right_transparency_texture[59][67] = 1;	doodle_right_transparency_texture[59][68] = 1;	doodle_right_transparency_texture[59][69] = 1;	doodle_right_transparency_texture[59][70] = 1;	doodle_right_transparency_texture[59][71] = 1;	doodle_right_transparency_texture[59][72] = 1;	doodle_right_transparency_texture[59][73] = 1;	doodle_right_transparency_texture[59][74] = 1;	doodle_right_transparency_texture[59][75] = 1;	doodle_right_transparency_texture[59][76] = 1;	doodle_right_transparency_texture[59][77] = 1;	doodle_right_transparency_texture[59][78] = 1;	doodle_right_transparency_texture[59][79] = 1;	doodle_right_transparency_texture[60][0] = 1;	doodle_right_transparency_texture[60][1] = 1;	doodle_right_transparency_texture[60][2] = 1;	doodle_right_transparency_texture[60][3] = 1;	doodle_right_transparency_texture[60][4] = 1;	doodle_right_transparency_texture[60][5] = 1;	doodle_right_transparency_texture[60][6] = 1;	doodle_right_transparency_texture[60][7] = 1;	doodle_right_transparency_texture[60][8] = 0;	doodle_right_transparency_texture[60][9] = 0;	doodle_right_transparency_texture[60][10] = 0;	doodle_right_transparency_texture[60][11] = 0;	doodle_right_transparency_texture[60][12] = 1;	doodle_right_transparency_texture[60][13] = 1;	doodle_right_transparency_texture[60][14] = 1;	doodle_right_transparency_texture[60][15] = 1;	doodle_right_transparency_texture[60][16] = 1;	doodle_right_transparency_texture[60][17] = 1;	doodle_right_transparency_texture[60][18] = 1;	doodle_right_transparency_texture[60][19] = 1;	doodle_right_transparency_texture[60][20] = 0;	doodle_right_transparency_texture[60][21] = 0;	doodle_right_transparency_texture[60][22] = 0;	doodle_right_transparency_texture[60][23] = 0;	doodle_right_transparency_texture[60][24] = 1;	doodle_right_transparency_texture[60][25] = 1;	doodle_right_transparency_texture[60][26] = 1;	doodle_right_transparency_texture[60][27] = 1;	doodle_right_transparency_texture[60][28] = 1;	doodle_right_transparency_texture[60][29] = 1;	doodle_right_transparency_texture[60][30] = 1;	doodle_right_transparency_texture[60][31] = 1;	doodle_right_transparency_texture[60][32] = 0;	doodle_right_transparency_texture[60][33] = 0;	doodle_right_transparency_texture[60][34] = 0;	doodle_right_transparency_texture[60][35] = 0;	doodle_right_transparency_texture[60][36] = 1;	doodle_right_transparency_texture[60][37] = 1;	doodle_right_transparency_texture[60][38] = 1;	doodle_right_transparency_texture[60][39] = 1;	doodle_right_transparency_texture[60][40] = 1;	doodle_right_transparency_texture[60][41] = 1;	doodle_right_transparency_texture[60][42] = 1;	doodle_right_transparency_texture[60][43] = 1;	doodle_right_transparency_texture[60][44] = 0;	doodle_right_transparency_texture[60][45] = 0;	doodle_right_transparency_texture[60][46] = 0;	doodle_right_transparency_texture[60][47] = 0;	doodle_right_transparency_texture[60][48] = 1;	doodle_right_transparency_texture[60][49] = 1;	doodle_right_transparency_texture[60][50] = 1;	doodle_right_transparency_texture[60][51] = 1;	doodle_right_transparency_texture[60][52] = 1;	doodle_right_transparency_texture[60][53] = 1;	doodle_right_transparency_texture[60][54] = 1;	doodle_right_transparency_texture[60][55] = 1;	doodle_right_transparency_texture[60][56] = 1;	doodle_right_transparency_texture[60][57] = 1;	doodle_right_transparency_texture[60][58] = 1;	doodle_right_transparency_texture[60][59] = 1;	doodle_right_transparency_texture[60][60] = 1;	doodle_right_transparency_texture[60][61] = 1;	doodle_right_transparency_texture[60][62] = 1;	doodle_right_transparency_texture[60][63] = 1;	doodle_right_transparency_texture[60][64] = 1;	doodle_right_transparency_texture[60][65] = 1;	doodle_right_transparency_texture[60][66] = 1;	doodle_right_transparency_texture[60][67] = 1;	doodle_right_transparency_texture[60][68] = 1;	doodle_right_transparency_texture[60][69] = 1;	doodle_right_transparency_texture[60][70] = 1;	doodle_right_transparency_texture[60][71] = 1;	doodle_right_transparency_texture[60][72] = 1;	doodle_right_transparency_texture[60][73] = 1;	doodle_right_transparency_texture[60][74] = 1;	doodle_right_transparency_texture[60][75] = 1;	doodle_right_transparency_texture[60][76] = 1;	doodle_right_transparency_texture[60][77] = 1;	doodle_right_transparency_texture[60][78] = 1;	doodle_right_transparency_texture[60][79] = 1;	doodle_right_transparency_texture[61][0] = 1;	doodle_right_transparency_texture[61][1] = 1;	doodle_right_transparency_texture[61][2] = 1;	doodle_right_transparency_texture[61][3] = 1;	doodle_right_transparency_texture[61][4] = 1;	doodle_right_transparency_texture[61][5] = 1;	doodle_right_transparency_texture[61][6] = 1;	doodle_right_transparency_texture[61][7] = 1;	doodle_right_transparency_texture[61][8] = 0;	doodle_right_transparency_texture[61][9] = 0;	doodle_right_transparency_texture[61][10] = 0;	doodle_right_transparency_texture[61][11] = 0;	doodle_right_transparency_texture[61][12] = 1;	doodle_right_transparency_texture[61][13] = 1;	doodle_right_transparency_texture[61][14] = 1;	doodle_right_transparency_texture[61][15] = 1;	doodle_right_transparency_texture[61][16] = 1;	doodle_right_transparency_texture[61][17] = 1;	doodle_right_transparency_texture[61][18] = 1;	doodle_right_transparency_texture[61][19] = 1;	doodle_right_transparency_texture[61][20] = 0;	doodle_right_transparency_texture[61][21] = 0;	doodle_right_transparency_texture[61][22] = 0;	doodle_right_transparency_texture[61][23] = 0;	doodle_right_transparency_texture[61][24] = 1;	doodle_right_transparency_texture[61][25] = 1;	doodle_right_transparency_texture[61][26] = 1;	doodle_right_transparency_texture[61][27] = 1;	doodle_right_transparency_texture[61][28] = 1;	doodle_right_transparency_texture[61][29] = 1;	doodle_right_transparency_texture[61][30] = 1;	doodle_right_transparency_texture[61][31] = 1;	doodle_right_transparency_texture[61][32] = 0;	doodle_right_transparency_texture[61][33] = 0;	doodle_right_transparency_texture[61][34] = 0;	doodle_right_transparency_texture[61][35] = 0;	doodle_right_transparency_texture[61][36] = 1;	doodle_right_transparency_texture[61][37] = 1;	doodle_right_transparency_texture[61][38] = 1;	doodle_right_transparency_texture[61][39] = 1;	doodle_right_transparency_texture[61][40] = 1;	doodle_right_transparency_texture[61][41] = 1;	doodle_right_transparency_texture[61][42] = 1;	doodle_right_transparency_texture[61][43] = 1;	doodle_right_transparency_texture[61][44] = 0;	doodle_right_transparency_texture[61][45] = 0;	doodle_right_transparency_texture[61][46] = 0;	doodle_right_transparency_texture[61][47] = 0;	doodle_right_transparency_texture[61][48] = 1;	doodle_right_transparency_texture[61][49] = 1;	doodle_right_transparency_texture[61][50] = 1;	doodle_right_transparency_texture[61][51] = 1;	doodle_right_transparency_texture[61][52] = 1;	doodle_right_transparency_texture[61][53] = 1;	doodle_right_transparency_texture[61][54] = 1;	doodle_right_transparency_texture[61][55] = 1;	doodle_right_transparency_texture[61][56] = 1;	doodle_right_transparency_texture[61][57] = 1;	doodle_right_transparency_texture[61][58] = 1;	doodle_right_transparency_texture[61][59] = 1;	doodle_right_transparency_texture[61][60] = 1;	doodle_right_transparency_texture[61][61] = 1;	doodle_right_transparency_texture[61][62] = 1;	doodle_right_transparency_texture[61][63] = 1;	doodle_right_transparency_texture[61][64] = 1;	doodle_right_transparency_texture[61][65] = 1;	doodle_right_transparency_texture[61][66] = 1;	doodle_right_transparency_texture[61][67] = 1;	doodle_right_transparency_texture[61][68] = 1;	doodle_right_transparency_texture[61][69] = 1;	doodle_right_transparency_texture[61][70] = 1;	doodle_right_transparency_texture[61][71] = 1;	doodle_right_transparency_texture[61][72] = 1;	doodle_right_transparency_texture[61][73] = 1;	doodle_right_transparency_texture[61][74] = 1;	doodle_right_transparency_texture[61][75] = 1;	doodle_right_transparency_texture[61][76] = 1;	doodle_right_transparency_texture[61][77] = 1;	doodle_right_transparency_texture[61][78] = 1;	doodle_right_transparency_texture[61][79] = 1;	doodle_right_transparency_texture[62][0] = 1;	doodle_right_transparency_texture[62][1] = 1;	doodle_right_transparency_texture[62][2] = 1;	doodle_right_transparency_texture[62][3] = 1;	doodle_right_transparency_texture[62][4] = 1;	doodle_right_transparency_texture[62][5] = 1;	doodle_right_transparency_texture[62][6] = 1;	doodle_right_transparency_texture[62][7] = 1;	doodle_right_transparency_texture[62][8] = 0;	doodle_right_transparency_texture[62][9] = 0;	doodle_right_transparency_texture[62][10] = 0;	doodle_right_transparency_texture[62][11] = 0;	doodle_right_transparency_texture[62][12] = 1;	doodle_right_transparency_texture[62][13] = 1;	doodle_right_transparency_texture[62][14] = 1;	doodle_right_transparency_texture[62][15] = 1;	doodle_right_transparency_texture[62][16] = 1;	doodle_right_transparency_texture[62][17] = 1;	doodle_right_transparency_texture[62][18] = 1;	doodle_right_transparency_texture[62][19] = 1;	doodle_right_transparency_texture[62][20] = 0;	doodle_right_transparency_texture[62][21] = 0;	doodle_right_transparency_texture[62][22] = 0;	doodle_right_transparency_texture[62][23] = 0;	doodle_right_transparency_texture[62][24] = 1;	doodle_right_transparency_texture[62][25] = 1;	doodle_right_transparency_texture[62][26] = 1;	doodle_right_transparency_texture[62][27] = 1;	doodle_right_transparency_texture[62][28] = 1;	doodle_right_transparency_texture[62][29] = 1;	doodle_right_transparency_texture[62][30] = 1;	doodle_right_transparency_texture[62][31] = 1;	doodle_right_transparency_texture[62][32] = 0;	doodle_right_transparency_texture[62][33] = 0;	doodle_right_transparency_texture[62][34] = 0;	doodle_right_transparency_texture[62][35] = 0;	doodle_right_transparency_texture[62][36] = 1;	doodle_right_transparency_texture[62][37] = 1;	doodle_right_transparency_texture[62][38] = 1;	doodle_right_transparency_texture[62][39] = 1;	doodle_right_transparency_texture[62][40] = 1;	doodle_right_transparency_texture[62][41] = 1;	doodle_right_transparency_texture[62][42] = 1;	doodle_right_transparency_texture[62][43] = 1;	doodle_right_transparency_texture[62][44] = 0;	doodle_right_transparency_texture[62][45] = 0;	doodle_right_transparency_texture[62][46] = 0;	doodle_right_transparency_texture[62][47] = 0;	doodle_right_transparency_texture[62][48] = 1;	doodle_right_transparency_texture[62][49] = 1;	doodle_right_transparency_texture[62][50] = 1;	doodle_right_transparency_texture[62][51] = 1;	doodle_right_transparency_texture[62][52] = 1;	doodle_right_transparency_texture[62][53] = 1;	doodle_right_transparency_texture[62][54] = 1;	doodle_right_transparency_texture[62][55] = 1;	doodle_right_transparency_texture[62][56] = 1;	doodle_right_transparency_texture[62][57] = 1;	doodle_right_transparency_texture[62][58] = 1;	doodle_right_transparency_texture[62][59] = 1;	doodle_right_transparency_texture[62][60] = 1;	doodle_right_transparency_texture[62][61] = 1;	doodle_right_transparency_texture[62][62] = 1;	doodle_right_transparency_texture[62][63] = 1;	doodle_right_transparency_texture[62][64] = 1;	doodle_right_transparency_texture[62][65] = 1;	doodle_right_transparency_texture[62][66] = 1;	doodle_right_transparency_texture[62][67] = 1;	doodle_right_transparency_texture[62][68] = 1;	doodle_right_transparency_texture[62][69] = 1;	doodle_right_transparency_texture[62][70] = 1;	doodle_right_transparency_texture[62][71] = 1;	doodle_right_transparency_texture[62][72] = 1;	doodle_right_transparency_texture[62][73] = 1;	doodle_right_transparency_texture[62][74] = 1;	doodle_right_transparency_texture[62][75] = 1;	doodle_right_transparency_texture[62][76] = 1;	doodle_right_transparency_texture[62][77] = 1;	doodle_right_transparency_texture[62][78] = 1;	doodle_right_transparency_texture[62][79] = 1;	doodle_right_transparency_texture[63][0] = 1;	doodle_right_transparency_texture[63][1] = 1;	doodle_right_transparency_texture[63][2] = 1;	doodle_right_transparency_texture[63][3] = 1;	doodle_right_transparency_texture[63][4] = 1;	doodle_right_transparency_texture[63][5] = 1;	doodle_right_transparency_texture[63][6] = 1;	doodle_right_transparency_texture[63][7] = 1;	doodle_right_transparency_texture[63][8] = 0;	doodle_right_transparency_texture[63][9] = 0;	doodle_right_transparency_texture[63][10] = 0;	doodle_right_transparency_texture[63][11] = 0;	doodle_right_transparency_texture[63][12] = 1;	doodle_right_transparency_texture[63][13] = 1;	doodle_right_transparency_texture[63][14] = 1;	doodle_right_transparency_texture[63][15] = 1;	doodle_right_transparency_texture[63][16] = 1;	doodle_right_transparency_texture[63][17] = 1;	doodle_right_transparency_texture[63][18] = 1;	doodle_right_transparency_texture[63][19] = 1;	doodle_right_transparency_texture[63][20] = 0;	doodle_right_transparency_texture[63][21] = 0;	doodle_right_transparency_texture[63][22] = 0;	doodle_right_transparency_texture[63][23] = 0;	doodle_right_transparency_texture[63][24] = 1;	doodle_right_transparency_texture[63][25] = 1;	doodle_right_transparency_texture[63][26] = 1;	doodle_right_transparency_texture[63][27] = 1;	doodle_right_transparency_texture[63][28] = 1;	doodle_right_transparency_texture[63][29] = 1;	doodle_right_transparency_texture[63][30] = 1;	doodle_right_transparency_texture[63][31] = 1;	doodle_right_transparency_texture[63][32] = 0;	doodle_right_transparency_texture[63][33] = 0;	doodle_right_transparency_texture[63][34] = 0;	doodle_right_transparency_texture[63][35] = 0;	doodle_right_transparency_texture[63][36] = 1;	doodle_right_transparency_texture[63][37] = 1;	doodle_right_transparency_texture[63][38] = 1;	doodle_right_transparency_texture[63][39] = 1;	doodle_right_transparency_texture[63][40] = 1;	doodle_right_transparency_texture[63][41] = 1;	doodle_right_transparency_texture[63][42] = 1;	doodle_right_transparency_texture[63][43] = 1;	doodle_right_transparency_texture[63][44] = 0;	doodle_right_transparency_texture[63][45] = 0;	doodle_right_transparency_texture[63][46] = 0;	doodle_right_transparency_texture[63][47] = 0;	doodle_right_transparency_texture[63][48] = 1;	doodle_right_transparency_texture[63][49] = 1;	doodle_right_transparency_texture[63][50] = 1;	doodle_right_transparency_texture[63][51] = 1;	doodle_right_transparency_texture[63][52] = 1;	doodle_right_transparency_texture[63][53] = 1;	doodle_right_transparency_texture[63][54] = 1;	doodle_right_transparency_texture[63][55] = 1;	doodle_right_transparency_texture[63][56] = 1;	doodle_right_transparency_texture[63][57] = 1;	doodle_right_transparency_texture[63][58] = 1;	doodle_right_transparency_texture[63][59] = 1;	doodle_right_transparency_texture[63][60] = 1;	doodle_right_transparency_texture[63][61] = 1;	doodle_right_transparency_texture[63][62] = 1;	doodle_right_transparency_texture[63][63] = 1;	doodle_right_transparency_texture[63][64] = 1;	doodle_right_transparency_texture[63][65] = 1;	doodle_right_transparency_texture[63][66] = 1;	doodle_right_transparency_texture[63][67] = 1;	doodle_right_transparency_texture[63][68] = 1;	doodle_right_transparency_texture[63][69] = 1;	doodle_right_transparency_texture[63][70] = 1;	doodle_right_transparency_texture[63][71] = 1;	doodle_right_transparency_texture[63][72] = 1;	doodle_right_transparency_texture[63][73] = 1;	doodle_right_transparency_texture[63][74] = 1;	doodle_right_transparency_texture[63][75] = 1;	doodle_right_transparency_texture[63][76] = 1;	doodle_right_transparency_texture[63][77] = 1;	doodle_right_transparency_texture[63][78] = 1;	doodle_right_transparency_texture[63][79] = 1;	doodle_right_transparency_texture[64][0] = 1;	doodle_right_transparency_texture[64][1] = 1;	doodle_right_transparency_texture[64][2] = 1;	doodle_right_transparency_texture[64][3] = 1;	doodle_right_transparency_texture[64][4] = 1;	doodle_right_transparency_texture[64][5] = 1;	doodle_right_transparency_texture[64][6] = 1;	doodle_right_transparency_texture[64][7] = 1;	doodle_right_transparency_texture[64][8] = 0;	doodle_right_transparency_texture[64][9] = 0;	doodle_right_transparency_texture[64][10] = 0;	doodle_right_transparency_texture[64][11] = 0;	doodle_right_transparency_texture[64][12] = 1;	doodle_right_transparency_texture[64][13] = 1;	doodle_right_transparency_texture[64][14] = 1;	doodle_right_transparency_texture[64][15] = 1;	doodle_right_transparency_texture[64][16] = 1;	doodle_right_transparency_texture[64][17] = 1;	doodle_right_transparency_texture[64][18] = 1;	doodle_right_transparency_texture[64][19] = 1;	doodle_right_transparency_texture[64][20] = 0;	doodle_right_transparency_texture[64][21] = 0;	doodle_right_transparency_texture[64][22] = 0;	doodle_right_transparency_texture[64][23] = 0;	doodle_right_transparency_texture[64][24] = 1;	doodle_right_transparency_texture[64][25] = 1;	doodle_right_transparency_texture[64][26] = 1;	doodle_right_transparency_texture[64][27] = 1;	doodle_right_transparency_texture[64][28] = 1;	doodle_right_transparency_texture[64][29] = 1;	doodle_right_transparency_texture[64][30] = 1;	doodle_right_transparency_texture[64][31] = 1;	doodle_right_transparency_texture[64][32] = 0;	doodle_right_transparency_texture[64][33] = 0;	doodle_right_transparency_texture[64][34] = 0;	doodle_right_transparency_texture[64][35] = 0;	doodle_right_transparency_texture[64][36] = 1;	doodle_right_transparency_texture[64][37] = 1;	doodle_right_transparency_texture[64][38] = 1;	doodle_right_transparency_texture[64][39] = 1;	doodle_right_transparency_texture[64][40] = 1;	doodle_right_transparency_texture[64][41] = 1;	doodle_right_transparency_texture[64][42] = 1;	doodle_right_transparency_texture[64][43] = 1;	doodle_right_transparency_texture[64][44] = 0;	doodle_right_transparency_texture[64][45] = 0;	doodle_right_transparency_texture[64][46] = 0;	doodle_right_transparency_texture[64][47] = 0;	doodle_right_transparency_texture[64][48] = 1;	doodle_right_transparency_texture[64][49] = 1;	doodle_right_transparency_texture[64][50] = 1;	doodle_right_transparency_texture[64][51] = 1;	doodle_right_transparency_texture[64][52] = 1;	doodle_right_transparency_texture[64][53] = 1;	doodle_right_transparency_texture[64][54] = 1;	doodle_right_transparency_texture[64][55] = 1;	doodle_right_transparency_texture[64][56] = 1;	doodle_right_transparency_texture[64][57] = 1;	doodle_right_transparency_texture[64][58] = 1;	doodle_right_transparency_texture[64][59] = 1;	doodle_right_transparency_texture[64][60] = 1;	doodle_right_transparency_texture[64][61] = 1;	doodle_right_transparency_texture[64][62] = 1;	doodle_right_transparency_texture[64][63] = 1;	doodle_right_transparency_texture[64][64] = 1;	doodle_right_transparency_texture[64][65] = 1;	doodle_right_transparency_texture[64][66] = 1;	doodle_right_transparency_texture[64][67] = 1;	doodle_right_transparency_texture[64][68] = 1;	doodle_right_transparency_texture[64][69] = 1;	doodle_right_transparency_texture[64][70] = 1;	doodle_right_transparency_texture[64][71] = 1;	doodle_right_transparency_texture[64][72] = 1;	doodle_right_transparency_texture[64][73] = 1;	doodle_right_transparency_texture[64][74] = 1;	doodle_right_transparency_texture[64][75] = 1;	doodle_right_transparency_texture[64][76] = 1;	doodle_right_transparency_texture[64][77] = 1;	doodle_right_transparency_texture[64][78] = 1;	doodle_right_transparency_texture[64][79] = 1;	doodle_right_transparency_texture[65][0] = 1;	doodle_right_transparency_texture[65][1] = 1;	doodle_right_transparency_texture[65][2] = 1;	doodle_right_transparency_texture[65][3] = 1;	doodle_right_transparency_texture[65][4] = 1;	doodle_right_transparency_texture[65][5] = 1;	doodle_right_transparency_texture[65][6] = 1;	doodle_right_transparency_texture[65][7] = 1;	doodle_right_transparency_texture[65][8] = 0;	doodle_right_transparency_texture[65][9] = 0;	doodle_right_transparency_texture[65][10] = 0;	doodle_right_transparency_texture[65][11] = 0;	doodle_right_transparency_texture[65][12] = 1;	doodle_right_transparency_texture[65][13] = 1;	doodle_right_transparency_texture[65][14] = 1;	doodle_right_transparency_texture[65][15] = 1;	doodle_right_transparency_texture[65][16] = 1;	doodle_right_transparency_texture[65][17] = 1;	doodle_right_transparency_texture[65][18] = 1;	doodle_right_transparency_texture[65][19] = 1;	doodle_right_transparency_texture[65][20] = 0;	doodle_right_transparency_texture[65][21] = 0;	doodle_right_transparency_texture[65][22] = 0;	doodle_right_transparency_texture[65][23] = 0;	doodle_right_transparency_texture[65][24] = 1;	doodle_right_transparency_texture[65][25] = 1;	doodle_right_transparency_texture[65][26] = 1;	doodle_right_transparency_texture[65][27] = 1;	doodle_right_transparency_texture[65][28] = 1;	doodle_right_transparency_texture[65][29] = 1;	doodle_right_transparency_texture[65][30] = 1;	doodle_right_transparency_texture[65][31] = 1;	doodle_right_transparency_texture[65][32] = 0;	doodle_right_transparency_texture[65][33] = 0;	doodle_right_transparency_texture[65][34] = 0;	doodle_right_transparency_texture[65][35] = 0;	doodle_right_transparency_texture[65][36] = 1;	doodle_right_transparency_texture[65][37] = 1;	doodle_right_transparency_texture[65][38] = 1;	doodle_right_transparency_texture[65][39] = 1;	doodle_right_transparency_texture[65][40] = 1;	doodle_right_transparency_texture[65][41] = 1;	doodle_right_transparency_texture[65][42] = 1;	doodle_right_transparency_texture[65][43] = 1;	doodle_right_transparency_texture[65][44] = 0;	doodle_right_transparency_texture[65][45] = 0;	doodle_right_transparency_texture[65][46] = 0;	doodle_right_transparency_texture[65][47] = 0;	doodle_right_transparency_texture[65][48] = 1;	doodle_right_transparency_texture[65][49] = 1;	doodle_right_transparency_texture[65][50] = 1;	doodle_right_transparency_texture[65][51] = 1;	doodle_right_transparency_texture[65][52] = 1;	doodle_right_transparency_texture[65][53] = 1;	doodle_right_transparency_texture[65][54] = 1;	doodle_right_transparency_texture[65][55] = 1;	doodle_right_transparency_texture[65][56] = 1;	doodle_right_transparency_texture[65][57] = 1;	doodle_right_transparency_texture[65][58] = 1;	doodle_right_transparency_texture[65][59] = 1;	doodle_right_transparency_texture[65][60] = 1;	doodle_right_transparency_texture[65][61] = 1;	doodle_right_transparency_texture[65][62] = 1;	doodle_right_transparency_texture[65][63] = 1;	doodle_right_transparency_texture[65][64] = 1;	doodle_right_transparency_texture[65][65] = 1;	doodle_right_transparency_texture[65][66] = 1;	doodle_right_transparency_texture[65][67] = 1;	doodle_right_transparency_texture[65][68] = 1;	doodle_right_transparency_texture[65][69] = 1;	doodle_right_transparency_texture[65][70] = 1;	doodle_right_transparency_texture[65][71] = 1;	doodle_right_transparency_texture[65][72] = 1;	doodle_right_transparency_texture[65][73] = 1;	doodle_right_transparency_texture[65][74] = 1;	doodle_right_transparency_texture[65][75] = 1;	doodle_right_transparency_texture[65][76] = 1;	doodle_right_transparency_texture[65][77] = 1;	doodle_right_transparency_texture[65][78] = 1;	doodle_right_transparency_texture[65][79] = 1;	doodle_right_transparency_texture[66][0] = 1;	doodle_right_transparency_texture[66][1] = 1;	doodle_right_transparency_texture[66][2] = 1;	doodle_right_transparency_texture[66][3] = 1;	doodle_right_transparency_texture[66][4] = 1;	doodle_right_transparency_texture[66][5] = 1;	doodle_right_transparency_texture[66][6] = 1;	doodle_right_transparency_texture[66][7] = 1;	doodle_right_transparency_texture[66][8] = 0;	doodle_right_transparency_texture[66][9] = 0;	doodle_right_transparency_texture[66][10] = 0;	doodle_right_transparency_texture[66][11] = 0;	doodle_right_transparency_texture[66][12] = 1;	doodle_right_transparency_texture[66][13] = 1;	doodle_right_transparency_texture[66][14] = 1;	doodle_right_transparency_texture[66][15] = 1;	doodle_right_transparency_texture[66][16] = 1;	doodle_right_transparency_texture[66][17] = 1;	doodle_right_transparency_texture[66][18] = 1;	doodle_right_transparency_texture[66][19] = 1;	doodle_right_transparency_texture[66][20] = 0;	doodle_right_transparency_texture[66][21] = 0;	doodle_right_transparency_texture[66][22] = 0;	doodle_right_transparency_texture[66][23] = 0;	doodle_right_transparency_texture[66][24] = 1;	doodle_right_transparency_texture[66][25] = 1;	doodle_right_transparency_texture[66][26] = 1;	doodle_right_transparency_texture[66][27] = 1;	doodle_right_transparency_texture[66][28] = 1;	doodle_right_transparency_texture[66][29] = 1;	doodle_right_transparency_texture[66][30] = 1;	doodle_right_transparency_texture[66][31] = 1;	doodle_right_transparency_texture[66][32] = 0;	doodle_right_transparency_texture[66][33] = 0;	doodle_right_transparency_texture[66][34] = 0;	doodle_right_transparency_texture[66][35] = 0;	doodle_right_transparency_texture[66][36] = 1;	doodle_right_transparency_texture[66][37] = 1;	doodle_right_transparency_texture[66][38] = 1;	doodle_right_transparency_texture[66][39] = 1;	doodle_right_transparency_texture[66][40] = 1;	doodle_right_transparency_texture[66][41] = 1;	doodle_right_transparency_texture[66][42] = 1;	doodle_right_transparency_texture[66][43] = 1;	doodle_right_transparency_texture[66][44] = 0;	doodle_right_transparency_texture[66][45] = 0;	doodle_right_transparency_texture[66][46] = 0;	doodle_right_transparency_texture[66][47] = 0;	doodle_right_transparency_texture[66][48] = 1;	doodle_right_transparency_texture[66][49] = 1;	doodle_right_transparency_texture[66][50] = 1;	doodle_right_transparency_texture[66][51] = 1;	doodle_right_transparency_texture[66][52] = 1;	doodle_right_transparency_texture[66][53] = 1;	doodle_right_transparency_texture[66][54] = 1;	doodle_right_transparency_texture[66][55] = 1;	doodle_right_transparency_texture[66][56] = 1;	doodle_right_transparency_texture[66][57] = 1;	doodle_right_transparency_texture[66][58] = 1;	doodle_right_transparency_texture[66][59] = 1;	doodle_right_transparency_texture[66][60] = 1;	doodle_right_transparency_texture[66][61] = 1;	doodle_right_transparency_texture[66][62] = 1;	doodle_right_transparency_texture[66][63] = 1;	doodle_right_transparency_texture[66][64] = 1;	doodle_right_transparency_texture[66][65] = 1;	doodle_right_transparency_texture[66][66] = 1;	doodle_right_transparency_texture[66][67] = 1;	doodle_right_transparency_texture[66][68] = 1;	doodle_right_transparency_texture[66][69] = 1;	doodle_right_transparency_texture[66][70] = 1;	doodle_right_transparency_texture[66][71] = 1;	doodle_right_transparency_texture[66][72] = 1;	doodle_right_transparency_texture[66][73] = 1;	doodle_right_transparency_texture[66][74] = 1;	doodle_right_transparency_texture[66][75] = 1;	doodle_right_transparency_texture[66][76] = 1;	doodle_right_transparency_texture[66][77] = 1;	doodle_right_transparency_texture[66][78] = 1;	doodle_right_transparency_texture[66][79] = 1;	doodle_right_transparency_texture[67][0] = 1;	doodle_right_transparency_texture[67][1] = 1;	doodle_right_transparency_texture[67][2] = 1;	doodle_right_transparency_texture[67][3] = 1;	doodle_right_transparency_texture[67][4] = 1;	doodle_right_transparency_texture[67][5] = 1;	doodle_right_transparency_texture[67][6] = 1;	doodle_right_transparency_texture[67][7] = 1;	doodle_right_transparency_texture[67][8] = 0;	doodle_right_transparency_texture[67][9] = 0;	doodle_right_transparency_texture[67][10] = 0;	doodle_right_transparency_texture[67][11] = 0;	doodle_right_transparency_texture[67][12] = 1;	doodle_right_transparency_texture[67][13] = 1;	doodle_right_transparency_texture[67][14] = 1;	doodle_right_transparency_texture[67][15] = 1;	doodle_right_transparency_texture[67][16] = 1;	doodle_right_transparency_texture[67][17] = 1;	doodle_right_transparency_texture[67][18] = 1;	doodle_right_transparency_texture[67][19] = 1;	doodle_right_transparency_texture[67][20] = 0;	doodle_right_transparency_texture[67][21] = 0;	doodle_right_transparency_texture[67][22] = 0;	doodle_right_transparency_texture[67][23] = 0;	doodle_right_transparency_texture[67][24] = 1;	doodle_right_transparency_texture[67][25] = 1;	doodle_right_transparency_texture[67][26] = 1;	doodle_right_transparency_texture[67][27] = 1;	doodle_right_transparency_texture[67][28] = 1;	doodle_right_transparency_texture[67][29] = 1;	doodle_right_transparency_texture[67][30] = 1;	doodle_right_transparency_texture[67][31] = 1;	doodle_right_transparency_texture[67][32] = 0;	doodle_right_transparency_texture[67][33] = 0;	doodle_right_transparency_texture[67][34] = 0;	doodle_right_transparency_texture[67][35] = 0;	doodle_right_transparency_texture[67][36] = 1;	doodle_right_transparency_texture[67][37] = 1;	doodle_right_transparency_texture[67][38] = 1;	doodle_right_transparency_texture[67][39] = 1;	doodle_right_transparency_texture[67][40] = 1;	doodle_right_transparency_texture[67][41] = 1;	doodle_right_transparency_texture[67][42] = 1;	doodle_right_transparency_texture[67][43] = 1;	doodle_right_transparency_texture[67][44] = 0;	doodle_right_transparency_texture[67][45] = 0;	doodle_right_transparency_texture[67][46] = 0;	doodle_right_transparency_texture[67][47] = 0;	doodle_right_transparency_texture[67][48] = 1;	doodle_right_transparency_texture[67][49] = 1;	doodle_right_transparency_texture[67][50] = 1;	doodle_right_transparency_texture[67][51] = 1;	doodle_right_transparency_texture[67][52] = 1;	doodle_right_transparency_texture[67][53] = 1;	doodle_right_transparency_texture[67][54] = 1;	doodle_right_transparency_texture[67][55] = 1;	doodle_right_transparency_texture[67][56] = 1;	doodle_right_transparency_texture[67][57] = 1;	doodle_right_transparency_texture[67][58] = 1;	doodle_right_transparency_texture[67][59] = 1;	doodle_right_transparency_texture[67][60] = 1;	doodle_right_transparency_texture[67][61] = 1;	doodle_right_transparency_texture[67][62] = 1;	doodle_right_transparency_texture[67][63] = 1;	doodle_right_transparency_texture[67][64] = 1;	doodle_right_transparency_texture[67][65] = 1;	doodle_right_transparency_texture[67][66] = 1;	doodle_right_transparency_texture[67][67] = 1;	doodle_right_transparency_texture[67][68] = 1;	doodle_right_transparency_texture[67][69] = 1;	doodle_right_transparency_texture[67][70] = 1;	doodle_right_transparency_texture[67][71] = 1;	doodle_right_transparency_texture[67][72] = 1;	doodle_right_transparency_texture[67][73] = 1;	doodle_right_transparency_texture[67][74] = 1;	doodle_right_transparency_texture[67][75] = 1;	doodle_right_transparency_texture[67][76] = 1;	doodle_right_transparency_texture[67][77] = 1;	doodle_right_transparency_texture[67][78] = 1;	doodle_right_transparency_texture[67][79] = 1;	doodle_right_transparency_texture[68][0] = 1;	doodle_right_transparency_texture[68][1] = 1;	doodle_right_transparency_texture[68][2] = 1;	doodle_right_transparency_texture[68][3] = 1;	doodle_right_transparency_texture[68][4] = 1;	doodle_right_transparency_texture[68][5] = 1;	doodle_right_transparency_texture[68][6] = 1;	doodle_right_transparency_texture[68][7] = 1;	doodle_right_transparency_texture[68][8] = 0;	doodle_right_transparency_texture[68][9] = 0;	doodle_right_transparency_texture[68][10] = 0;	doodle_right_transparency_texture[68][11] = 0;	doodle_right_transparency_texture[68][12] = 0;	doodle_right_transparency_texture[68][13] = 0;	doodle_right_transparency_texture[68][14] = 0;	doodle_right_transparency_texture[68][15] = 0;	doodle_right_transparency_texture[68][16] = 1;	doodle_right_transparency_texture[68][17] = 1;	doodle_right_transparency_texture[68][18] = 1;	doodle_right_transparency_texture[68][19] = 1;	doodle_right_transparency_texture[68][20] = 0;	doodle_right_transparency_texture[68][21] = 0;	doodle_right_transparency_texture[68][22] = 0;	doodle_right_transparency_texture[68][23] = 0;	doodle_right_transparency_texture[68][24] = 0;	doodle_right_transparency_texture[68][25] = 0;	doodle_right_transparency_texture[68][26] = 0;	doodle_right_transparency_texture[68][27] = 0;	doodle_right_transparency_texture[68][28] = 1;	doodle_right_transparency_texture[68][29] = 1;	doodle_right_transparency_texture[68][30] = 1;	doodle_right_transparency_texture[68][31] = 1;	doodle_right_transparency_texture[68][32] = 0;	doodle_right_transparency_texture[68][33] = 0;	doodle_right_transparency_texture[68][34] = 0;	doodle_right_transparency_texture[68][35] = 0;	doodle_right_transparency_texture[68][36] = 0;	doodle_right_transparency_texture[68][37] = 0;	doodle_right_transparency_texture[68][38] = 0;	doodle_right_transparency_texture[68][39] = 0;	doodle_right_transparency_texture[68][40] = 1;	doodle_right_transparency_texture[68][41] = 1;	doodle_right_transparency_texture[68][42] = 1;	doodle_right_transparency_texture[68][43] = 1;	doodle_right_transparency_texture[68][44] = 0;	doodle_right_transparency_texture[68][45] = 0;	doodle_right_transparency_texture[68][46] = 0;	doodle_right_transparency_texture[68][47] = 0;	doodle_right_transparency_texture[68][48] = 0;	doodle_right_transparency_texture[68][49] = 0;	doodle_right_transparency_texture[68][50] = 0;	doodle_right_transparency_texture[68][51] = 0;	doodle_right_transparency_texture[68][52] = 1;	doodle_right_transparency_texture[68][53] = 1;	doodle_right_transparency_texture[68][54] = 1;	doodle_right_transparency_texture[68][55] = 1;	doodle_right_transparency_texture[68][56] = 1;	doodle_right_transparency_texture[68][57] = 1;	doodle_right_transparency_texture[68][58] = 1;	doodle_right_transparency_texture[68][59] = 1;	doodle_right_transparency_texture[68][60] = 1;	doodle_right_transparency_texture[68][61] = 1;	doodle_right_transparency_texture[68][62] = 1;	doodle_right_transparency_texture[68][63] = 1;	doodle_right_transparency_texture[68][64] = 1;	doodle_right_transparency_texture[68][65] = 1;	doodle_right_transparency_texture[68][66] = 1;	doodle_right_transparency_texture[68][67] = 1;	doodle_right_transparency_texture[68][68] = 1;	doodle_right_transparency_texture[68][69] = 1;	doodle_right_transparency_texture[68][70] = 1;	doodle_right_transparency_texture[68][71] = 1;	doodle_right_transparency_texture[68][72] = 1;	doodle_right_transparency_texture[68][73] = 1;	doodle_right_transparency_texture[68][74] = 1;	doodle_right_transparency_texture[68][75] = 1;	doodle_right_transparency_texture[68][76] = 1;	doodle_right_transparency_texture[68][77] = 1;	doodle_right_transparency_texture[68][78] = 1;	doodle_right_transparency_texture[68][79] = 1;	doodle_right_transparency_texture[69][0] = 1;	doodle_right_transparency_texture[69][1] = 1;	doodle_right_transparency_texture[69][2] = 1;	doodle_right_transparency_texture[69][3] = 1;	doodle_right_transparency_texture[69][4] = 1;	doodle_right_transparency_texture[69][5] = 1;	doodle_right_transparency_texture[69][6] = 1;	doodle_right_transparency_texture[69][7] = 1;	doodle_right_transparency_texture[69][8] = 0;	doodle_right_transparency_texture[69][9] = 0;	doodle_right_transparency_texture[69][10] = 0;	doodle_right_transparency_texture[69][11] = 0;	doodle_right_transparency_texture[69][12] = 0;	doodle_right_transparency_texture[69][13] = 0;	doodle_right_transparency_texture[69][14] = 0;	doodle_right_transparency_texture[69][15] = 0;	doodle_right_transparency_texture[69][16] = 1;	doodle_right_transparency_texture[69][17] = 1;	doodle_right_transparency_texture[69][18] = 1;	doodle_right_transparency_texture[69][19] = 1;	doodle_right_transparency_texture[69][20] = 0;	doodle_right_transparency_texture[69][21] = 0;	doodle_right_transparency_texture[69][22] = 0;	doodle_right_transparency_texture[69][23] = 0;	doodle_right_transparency_texture[69][24] = 0;	doodle_right_transparency_texture[69][25] = 0;	doodle_right_transparency_texture[69][26] = 0;	doodle_right_transparency_texture[69][27] = 0;	doodle_right_transparency_texture[69][28] = 1;	doodle_right_transparency_texture[69][29] = 1;	doodle_right_transparency_texture[69][30] = 1;	doodle_right_transparency_texture[69][31] = 1;	doodle_right_transparency_texture[69][32] = 0;	doodle_right_transparency_texture[69][33] = 0;	doodle_right_transparency_texture[69][34] = 0;	doodle_right_transparency_texture[69][35] = 0;	doodle_right_transparency_texture[69][36] = 0;	doodle_right_transparency_texture[69][37] = 0;	doodle_right_transparency_texture[69][38] = 0;	doodle_right_transparency_texture[69][39] = 0;	doodle_right_transparency_texture[69][40] = 1;	doodle_right_transparency_texture[69][41] = 1;	doodle_right_transparency_texture[69][42] = 1;	doodle_right_transparency_texture[69][43] = 1;	doodle_right_transparency_texture[69][44] = 0;	doodle_right_transparency_texture[69][45] = 0;	doodle_right_transparency_texture[69][46] = 0;	doodle_right_transparency_texture[69][47] = 0;	doodle_right_transparency_texture[69][48] = 0;	doodle_right_transparency_texture[69][49] = 0;	doodle_right_transparency_texture[69][50] = 0;	doodle_right_transparency_texture[69][51] = 0;	doodle_right_transparency_texture[69][52] = 1;	doodle_right_transparency_texture[69][53] = 1;	doodle_right_transparency_texture[69][54] = 1;	doodle_right_transparency_texture[69][55] = 1;	doodle_right_transparency_texture[69][56] = 1;	doodle_right_transparency_texture[69][57] = 1;	doodle_right_transparency_texture[69][58] = 1;	doodle_right_transparency_texture[69][59] = 1;	doodle_right_transparency_texture[69][60] = 1;	doodle_right_transparency_texture[69][61] = 1;	doodle_right_transparency_texture[69][62] = 1;	doodle_right_transparency_texture[69][63] = 1;	doodle_right_transparency_texture[69][64] = 1;	doodle_right_transparency_texture[69][65] = 1;	doodle_right_transparency_texture[69][66] = 1;	doodle_right_transparency_texture[69][67] = 1;	doodle_right_transparency_texture[69][68] = 1;	doodle_right_transparency_texture[69][69] = 1;	doodle_right_transparency_texture[69][70] = 1;	doodle_right_transparency_texture[69][71] = 1;	doodle_right_transparency_texture[69][72] = 1;	doodle_right_transparency_texture[69][73] = 1;	doodle_right_transparency_texture[69][74] = 1;	doodle_right_transparency_texture[69][75] = 1;	doodle_right_transparency_texture[69][76] = 1;	doodle_right_transparency_texture[69][77] = 1;	doodle_right_transparency_texture[69][78] = 1;	doodle_right_transparency_texture[69][79] = 1;	doodle_right_transparency_texture[70][0] = 1;	doodle_right_transparency_texture[70][1] = 1;	doodle_right_transparency_texture[70][2] = 1;	doodle_right_transparency_texture[70][3] = 1;	doodle_right_transparency_texture[70][4] = 1;	doodle_right_transparency_texture[70][5] = 1;	doodle_right_transparency_texture[70][6] = 1;	doodle_right_transparency_texture[70][7] = 1;	doodle_right_transparency_texture[70][8] = 0;	doodle_right_transparency_texture[70][9] = 0;	doodle_right_transparency_texture[70][10] = 0;	doodle_right_transparency_texture[70][11] = 0;	doodle_right_transparency_texture[70][12] = 0;	doodle_right_transparency_texture[70][13] = 0;	doodle_right_transparency_texture[70][14] = 0;	doodle_right_transparency_texture[70][15] = 0;	doodle_right_transparency_texture[70][16] = 1;	doodle_right_transparency_texture[70][17] = 1;	doodle_right_transparency_texture[70][18] = 1;	doodle_right_transparency_texture[70][19] = 1;	doodle_right_transparency_texture[70][20] = 0;	doodle_right_transparency_texture[70][21] = 0;	doodle_right_transparency_texture[70][22] = 0;	doodle_right_transparency_texture[70][23] = 0;	doodle_right_transparency_texture[70][24] = 0;	doodle_right_transparency_texture[70][25] = 0;	doodle_right_transparency_texture[70][26] = 0;	doodle_right_transparency_texture[70][27] = 0;	doodle_right_transparency_texture[70][28] = 1;	doodle_right_transparency_texture[70][29] = 1;	doodle_right_transparency_texture[70][30] = 1;	doodle_right_transparency_texture[70][31] = 1;	doodle_right_transparency_texture[70][32] = 0;	doodle_right_transparency_texture[70][33] = 0;	doodle_right_transparency_texture[70][34] = 0;	doodle_right_transparency_texture[70][35] = 0;	doodle_right_transparency_texture[70][36] = 0;	doodle_right_transparency_texture[70][37] = 0;	doodle_right_transparency_texture[70][38] = 0;	doodle_right_transparency_texture[70][39] = 0;	doodle_right_transparency_texture[70][40] = 1;	doodle_right_transparency_texture[70][41] = 1;	doodle_right_transparency_texture[70][42] = 1;	doodle_right_transparency_texture[70][43] = 1;	doodle_right_transparency_texture[70][44] = 0;	doodle_right_transparency_texture[70][45] = 0;	doodle_right_transparency_texture[70][46] = 0;	doodle_right_transparency_texture[70][47] = 0;	doodle_right_transparency_texture[70][48] = 0;	doodle_right_transparency_texture[70][49] = 0;	doodle_right_transparency_texture[70][50] = 0;	doodle_right_transparency_texture[70][51] = 0;	doodle_right_transparency_texture[70][52] = 1;	doodle_right_transparency_texture[70][53] = 1;	doodle_right_transparency_texture[70][54] = 1;	doodle_right_transparency_texture[70][55] = 1;	doodle_right_transparency_texture[70][56] = 1;	doodle_right_transparency_texture[70][57] = 1;	doodle_right_transparency_texture[70][58] = 1;	doodle_right_transparency_texture[70][59] = 1;	doodle_right_transparency_texture[70][60] = 1;	doodle_right_transparency_texture[70][61] = 1;	doodle_right_transparency_texture[70][62] = 1;	doodle_right_transparency_texture[70][63] = 1;	doodle_right_transparency_texture[70][64] = 1;	doodle_right_transparency_texture[70][65] = 1;	doodle_right_transparency_texture[70][66] = 1;	doodle_right_transparency_texture[70][67] = 1;	doodle_right_transparency_texture[70][68] = 1;	doodle_right_transparency_texture[70][69] = 1;	doodle_right_transparency_texture[70][70] = 1;	doodle_right_transparency_texture[70][71] = 1;	doodle_right_transparency_texture[70][72] = 1;	doodle_right_transparency_texture[70][73] = 1;	doodle_right_transparency_texture[70][74] = 1;	doodle_right_transparency_texture[70][75] = 1;	doodle_right_transparency_texture[70][76] = 1;	doodle_right_transparency_texture[70][77] = 1;	doodle_right_transparency_texture[70][78] = 1;	doodle_right_transparency_texture[70][79] = 1;	doodle_right_transparency_texture[71][0] = 1;	doodle_right_transparency_texture[71][1] = 1;	doodle_right_transparency_texture[71][2] = 1;	doodle_right_transparency_texture[71][3] = 1;	doodle_right_transparency_texture[71][4] = 1;	doodle_right_transparency_texture[71][5] = 1;	doodle_right_transparency_texture[71][6] = 1;	doodle_right_transparency_texture[71][7] = 1;	doodle_right_transparency_texture[71][8] = 0;	doodle_right_transparency_texture[71][9] = 0;	doodle_right_transparency_texture[71][10] = 0;	doodle_right_transparency_texture[71][11] = 0;	doodle_right_transparency_texture[71][12] = 0;	doodle_right_transparency_texture[71][13] = 0;	doodle_right_transparency_texture[71][14] = 0;	doodle_right_transparency_texture[71][15] = 0;	doodle_right_transparency_texture[71][16] = 1;	doodle_right_transparency_texture[71][17] = 1;	doodle_right_transparency_texture[71][18] = 1;	doodle_right_transparency_texture[71][19] = 1;	doodle_right_transparency_texture[71][20] = 0;	doodle_right_transparency_texture[71][21] = 0;	doodle_right_transparency_texture[71][22] = 0;	doodle_right_transparency_texture[71][23] = 0;	doodle_right_transparency_texture[71][24] = 0;	doodle_right_transparency_texture[71][25] = 0;	doodle_right_transparency_texture[71][26] = 0;	doodle_right_transparency_texture[71][27] = 0;	doodle_right_transparency_texture[71][28] = 1;	doodle_right_transparency_texture[71][29] = 1;	doodle_right_transparency_texture[71][30] = 1;	doodle_right_transparency_texture[71][31] = 1;	doodle_right_transparency_texture[71][32] = 0;	doodle_right_transparency_texture[71][33] = 0;	doodle_right_transparency_texture[71][34] = 0;	doodle_right_transparency_texture[71][35] = 0;	doodle_right_transparency_texture[71][36] = 0;	doodle_right_transparency_texture[71][37] = 0;	doodle_right_transparency_texture[71][38] = 0;	doodle_right_transparency_texture[71][39] = 0;	doodle_right_transparency_texture[71][40] = 1;	doodle_right_transparency_texture[71][41] = 1;	doodle_right_transparency_texture[71][42] = 1;	doodle_right_transparency_texture[71][43] = 1;	doodle_right_transparency_texture[71][44] = 0;	doodle_right_transparency_texture[71][45] = 0;	doodle_right_transparency_texture[71][46] = 0;	doodle_right_transparency_texture[71][47] = 0;	doodle_right_transparency_texture[71][48] = 0;	doodle_right_transparency_texture[71][49] = 0;	doodle_right_transparency_texture[71][50] = 0;	doodle_right_transparency_texture[71][51] = 0;	doodle_right_transparency_texture[71][52] = 1;	doodle_right_transparency_texture[71][53] = 1;	doodle_right_transparency_texture[71][54] = 1;	doodle_right_transparency_texture[71][55] = 1;	doodle_right_transparency_texture[71][56] = 1;	doodle_right_transparency_texture[71][57] = 1;	doodle_right_transparency_texture[71][58] = 1;	doodle_right_transparency_texture[71][59] = 1;	doodle_right_transparency_texture[71][60] = 1;	doodle_right_transparency_texture[71][61] = 1;	doodle_right_transparency_texture[71][62] = 1;	doodle_right_transparency_texture[71][63] = 1;	doodle_right_transparency_texture[71][64] = 1;	doodle_right_transparency_texture[71][65] = 1;	doodle_right_transparency_texture[71][66] = 1;	doodle_right_transparency_texture[71][67] = 1;	doodle_right_transparency_texture[71][68] = 1;	doodle_right_transparency_texture[71][69] = 1;	doodle_right_transparency_texture[71][70] = 1;	doodle_right_transparency_texture[71][71] = 1;	doodle_right_transparency_texture[71][72] = 1;	doodle_right_transparency_texture[71][73] = 1;	doodle_right_transparency_texture[71][74] = 1;	doodle_right_transparency_texture[71][75] = 1;	doodle_right_transparency_texture[71][76] = 1;	doodle_right_transparency_texture[71][77] = 1;	doodle_right_transparency_texture[71][78] = 1;	doodle_right_transparency_texture[71][79] = 1;	doodle_right_transparency_texture[72][0] = 1;	doodle_right_transparency_texture[72][1] = 1;	doodle_right_transparency_texture[72][2] = 1;	doodle_right_transparency_texture[72][3] = 1;	doodle_right_transparency_texture[72][4] = 1;	doodle_right_transparency_texture[72][5] = 1;	doodle_right_transparency_texture[72][6] = 1;	doodle_right_transparency_texture[72][7] = 1;	doodle_right_transparency_texture[72][8] = 1;	doodle_right_transparency_texture[72][9] = 1;	doodle_right_transparency_texture[72][10] = 1;	doodle_right_transparency_texture[72][11] = 1;	doodle_right_transparency_texture[72][12] = 1;	doodle_right_transparency_texture[72][13] = 1;	doodle_right_transparency_texture[72][14] = 1;	doodle_right_transparency_texture[72][15] = 1;	doodle_right_transparency_texture[72][16] = 1;	doodle_right_transparency_texture[72][17] = 1;	doodle_right_transparency_texture[72][18] = 1;	doodle_right_transparency_texture[72][19] = 1;	doodle_right_transparency_texture[72][20] = 1;	doodle_right_transparency_texture[72][21] = 1;	doodle_right_transparency_texture[72][22] = 1;	doodle_right_transparency_texture[72][23] = 1;	doodle_right_transparency_texture[72][24] = 1;	doodle_right_transparency_texture[72][25] = 1;	doodle_right_transparency_texture[72][26] = 1;	doodle_right_transparency_texture[72][27] = 1;	doodle_right_transparency_texture[72][28] = 1;	doodle_right_transparency_texture[72][29] = 1;	doodle_right_transparency_texture[72][30] = 1;	doodle_right_transparency_texture[72][31] = 1;	doodle_right_transparency_texture[72][32] = 1;	doodle_right_transparency_texture[72][33] = 1;	doodle_right_transparency_texture[72][34] = 1;	doodle_right_transparency_texture[72][35] = 1;	doodle_right_transparency_texture[72][36] = 1;	doodle_right_transparency_texture[72][37] = 1;	doodle_right_transparency_texture[72][38] = 1;	doodle_right_transparency_texture[72][39] = 1;	doodle_right_transparency_texture[72][40] = 1;	doodle_right_transparency_texture[72][41] = 1;	doodle_right_transparency_texture[72][42] = 1;	doodle_right_transparency_texture[72][43] = 1;	doodle_right_transparency_texture[72][44] = 1;	doodle_right_transparency_texture[72][45] = 1;	doodle_right_transparency_texture[72][46] = 1;	doodle_right_transparency_texture[72][47] = 1;	doodle_right_transparency_texture[72][48] = 1;	doodle_right_transparency_texture[72][49] = 1;	doodle_right_transparency_texture[72][50] = 1;	doodle_right_transparency_texture[72][51] = 1;	doodle_right_transparency_texture[72][52] = 1;	doodle_right_transparency_texture[72][53] = 1;	doodle_right_transparency_texture[72][54] = 1;	doodle_right_transparency_texture[72][55] = 1;	doodle_right_transparency_texture[72][56] = 1;	doodle_right_transparency_texture[72][57] = 1;	doodle_right_transparency_texture[72][58] = 1;	doodle_right_transparency_texture[72][59] = 1;	doodle_right_transparency_texture[72][60] = 1;	doodle_right_transparency_texture[72][61] = 1;	doodle_right_transparency_texture[72][62] = 1;	doodle_right_transparency_texture[72][63] = 1;	doodle_right_transparency_texture[72][64] = 1;	doodle_right_transparency_texture[72][65] = 1;	doodle_right_transparency_texture[72][66] = 1;	doodle_right_transparency_texture[72][67] = 1;	doodle_right_transparency_texture[72][68] = 1;	doodle_right_transparency_texture[72][69] = 1;	doodle_right_transparency_texture[72][70] = 1;	doodle_right_transparency_texture[72][71] = 1;	doodle_right_transparency_texture[72][72] = 1;	doodle_right_transparency_texture[72][73] = 1;	doodle_right_transparency_texture[72][74] = 1;	doodle_right_transparency_texture[72][75] = 1;	doodle_right_transparency_texture[72][76] = 1;	doodle_right_transparency_texture[72][77] = 1;	doodle_right_transparency_texture[72][78] = 1;	doodle_right_transparency_texture[72][79] = 1;	doodle_right_transparency_texture[73][0] = 1;	doodle_right_transparency_texture[73][1] = 1;	doodle_right_transparency_texture[73][2] = 1;	doodle_right_transparency_texture[73][3] = 1;	doodle_right_transparency_texture[73][4] = 1;	doodle_right_transparency_texture[73][5] = 1;	doodle_right_transparency_texture[73][6] = 1;	doodle_right_transparency_texture[73][7] = 1;	doodle_right_transparency_texture[73][8] = 1;	doodle_right_transparency_texture[73][9] = 1;	doodle_right_transparency_texture[73][10] = 1;	doodle_right_transparency_texture[73][11] = 1;	doodle_right_transparency_texture[73][12] = 1;	doodle_right_transparency_texture[73][13] = 1;	doodle_right_transparency_texture[73][14] = 1;	doodle_right_transparency_texture[73][15] = 1;	doodle_right_transparency_texture[73][16] = 1;	doodle_right_transparency_texture[73][17] = 1;	doodle_right_transparency_texture[73][18] = 1;	doodle_right_transparency_texture[73][19] = 1;	doodle_right_transparency_texture[73][20] = 1;	doodle_right_transparency_texture[73][21] = 1;	doodle_right_transparency_texture[73][22] = 1;	doodle_right_transparency_texture[73][23] = 1;	doodle_right_transparency_texture[73][24] = 1;	doodle_right_transparency_texture[73][25] = 1;	doodle_right_transparency_texture[73][26] = 1;	doodle_right_transparency_texture[73][27] = 1;	doodle_right_transparency_texture[73][28] = 1;	doodle_right_transparency_texture[73][29] = 1;	doodle_right_transparency_texture[73][30] = 1;	doodle_right_transparency_texture[73][31] = 1;	doodle_right_transparency_texture[73][32] = 1;	doodle_right_transparency_texture[73][33] = 1;	doodle_right_transparency_texture[73][34] = 1;	doodle_right_transparency_texture[73][35] = 1;	doodle_right_transparency_texture[73][36] = 1;	doodle_right_transparency_texture[73][37] = 1;	doodle_right_transparency_texture[73][38] = 1;	doodle_right_transparency_texture[73][39] = 1;	doodle_right_transparency_texture[73][40] = 1;	doodle_right_transparency_texture[73][41] = 1;	doodle_right_transparency_texture[73][42] = 1;	doodle_right_transparency_texture[73][43] = 1;	doodle_right_transparency_texture[73][44] = 1;	doodle_right_transparency_texture[73][45] = 1;	doodle_right_transparency_texture[73][46] = 1;	doodle_right_transparency_texture[73][47] = 1;	doodle_right_transparency_texture[73][48] = 1;	doodle_right_transparency_texture[73][49] = 1;	doodle_right_transparency_texture[73][50] = 1;	doodle_right_transparency_texture[73][51] = 1;	doodle_right_transparency_texture[73][52] = 1;	doodle_right_transparency_texture[73][53] = 1;	doodle_right_transparency_texture[73][54] = 1;	doodle_right_transparency_texture[73][55] = 1;	doodle_right_transparency_texture[73][56] = 1;	doodle_right_transparency_texture[73][57] = 1;	doodle_right_transparency_texture[73][58] = 1;	doodle_right_transparency_texture[73][59] = 1;	doodle_right_transparency_texture[73][60] = 1;	doodle_right_transparency_texture[73][61] = 1;	doodle_right_transparency_texture[73][62] = 1;	doodle_right_transparency_texture[73][63] = 1;	doodle_right_transparency_texture[73][64] = 1;	doodle_right_transparency_texture[73][65] = 1;	doodle_right_transparency_texture[73][66] = 1;	doodle_right_transparency_texture[73][67] = 1;	doodle_right_transparency_texture[73][68] = 1;	doodle_right_transparency_texture[73][69] = 1;	doodle_right_transparency_texture[73][70] = 1;	doodle_right_transparency_texture[73][71] = 1;	doodle_right_transparency_texture[73][72] = 1;	doodle_right_transparency_texture[73][73] = 1;	doodle_right_transparency_texture[73][74] = 1;	doodle_right_transparency_texture[73][75] = 1;	doodle_right_transparency_texture[73][76] = 1;	doodle_right_transparency_texture[73][77] = 1;	doodle_right_transparency_texture[73][78] = 1;	doodle_right_transparency_texture[73][79] = 1;	doodle_right_transparency_texture[74][0] = 1;	doodle_right_transparency_texture[74][1] = 1;	doodle_right_transparency_texture[74][2] = 1;	doodle_right_transparency_texture[74][3] = 1;	doodle_right_transparency_texture[74][4] = 1;	doodle_right_transparency_texture[74][5] = 1;	doodle_right_transparency_texture[74][6] = 1;	doodle_right_transparency_texture[74][7] = 1;	doodle_right_transparency_texture[74][8] = 1;	doodle_right_transparency_texture[74][9] = 1;	doodle_right_transparency_texture[74][10] = 1;	doodle_right_transparency_texture[74][11] = 1;	doodle_right_transparency_texture[74][12] = 1;	doodle_right_transparency_texture[74][13] = 1;	doodle_right_transparency_texture[74][14] = 1;	doodle_right_transparency_texture[74][15] = 1;	doodle_right_transparency_texture[74][16] = 1;	doodle_right_transparency_texture[74][17] = 1;	doodle_right_transparency_texture[74][18] = 1;	doodle_right_transparency_texture[74][19] = 1;	doodle_right_transparency_texture[74][20] = 1;	doodle_right_transparency_texture[74][21] = 1;	doodle_right_transparency_texture[74][22] = 1;	doodle_right_transparency_texture[74][23] = 1;	doodle_right_transparency_texture[74][24] = 1;	doodle_right_transparency_texture[74][25] = 1;	doodle_right_transparency_texture[74][26] = 1;	doodle_right_transparency_texture[74][27] = 1;	doodle_right_transparency_texture[74][28] = 1;	doodle_right_transparency_texture[74][29] = 1;	doodle_right_transparency_texture[74][30] = 1;	doodle_right_transparency_texture[74][31] = 1;	doodle_right_transparency_texture[74][32] = 1;	doodle_right_transparency_texture[74][33] = 1;	doodle_right_transparency_texture[74][34] = 1;	doodle_right_transparency_texture[74][35] = 1;	doodle_right_transparency_texture[74][36] = 1;	doodle_right_transparency_texture[74][37] = 1;	doodle_right_transparency_texture[74][38] = 1;	doodle_right_transparency_texture[74][39] = 1;	doodle_right_transparency_texture[74][40] = 1;	doodle_right_transparency_texture[74][41] = 1;	doodle_right_transparency_texture[74][42] = 1;	doodle_right_transparency_texture[74][43] = 1;	doodle_right_transparency_texture[74][44] = 1;	doodle_right_transparency_texture[74][45] = 1;	doodle_right_transparency_texture[74][46] = 1;	doodle_right_transparency_texture[74][47] = 1;	doodle_right_transparency_texture[74][48] = 1;	doodle_right_transparency_texture[74][49] = 1;	doodle_right_transparency_texture[74][50] = 1;	doodle_right_transparency_texture[74][51] = 1;	doodle_right_transparency_texture[74][52] = 1;	doodle_right_transparency_texture[74][53] = 1;	doodle_right_transparency_texture[74][54] = 1;	doodle_right_transparency_texture[74][55] = 1;	doodle_right_transparency_texture[74][56] = 1;	doodle_right_transparency_texture[74][57] = 1;	doodle_right_transparency_texture[74][58] = 1;	doodle_right_transparency_texture[74][59] = 1;	doodle_right_transparency_texture[74][60] = 1;	doodle_right_transparency_texture[74][61] = 1;	doodle_right_transparency_texture[74][62] = 1;	doodle_right_transparency_texture[74][63] = 1;	doodle_right_transparency_texture[74][64] = 1;	doodle_right_transparency_texture[74][65] = 1;	doodle_right_transparency_texture[74][66] = 1;	doodle_right_transparency_texture[74][67] = 1;	doodle_right_transparency_texture[74][68] = 1;	doodle_right_transparency_texture[74][69] = 1;	doodle_right_transparency_texture[74][70] = 1;	doodle_right_transparency_texture[74][71] = 1;	doodle_right_transparency_texture[74][72] = 1;	doodle_right_transparency_texture[74][73] = 1;	doodle_right_transparency_texture[74][74] = 1;	doodle_right_transparency_texture[74][75] = 1;	doodle_right_transparency_texture[74][76] = 1;	doodle_right_transparency_texture[74][77] = 1;	doodle_right_transparency_texture[74][78] = 1;	doodle_right_transparency_texture[74][79] = 1;	doodle_right_transparency_texture[75][0] = 1;	doodle_right_transparency_texture[75][1] = 1;	doodle_right_transparency_texture[75][2] = 1;	doodle_right_transparency_texture[75][3] = 1;	doodle_right_transparency_texture[75][4] = 1;	doodle_right_transparency_texture[75][5] = 1;	doodle_right_transparency_texture[75][6] = 1;	doodle_right_transparency_texture[75][7] = 1;	doodle_right_transparency_texture[75][8] = 1;	doodle_right_transparency_texture[75][9] = 1;	doodle_right_transparency_texture[75][10] = 1;	doodle_right_transparency_texture[75][11] = 1;	doodle_right_transparency_texture[75][12] = 1;	doodle_right_transparency_texture[75][13] = 1;	doodle_right_transparency_texture[75][14] = 1;	doodle_right_transparency_texture[75][15] = 1;	doodle_right_transparency_texture[75][16] = 1;	doodle_right_transparency_texture[75][17] = 1;	doodle_right_transparency_texture[75][18] = 1;	doodle_right_transparency_texture[75][19] = 1;	doodle_right_transparency_texture[75][20] = 1;	doodle_right_transparency_texture[75][21] = 1;	doodle_right_transparency_texture[75][22] = 1;	doodle_right_transparency_texture[75][23] = 1;	doodle_right_transparency_texture[75][24] = 1;	doodle_right_transparency_texture[75][25] = 1;	doodle_right_transparency_texture[75][26] = 1;	doodle_right_transparency_texture[75][27] = 1;	doodle_right_transparency_texture[75][28] = 1;	doodle_right_transparency_texture[75][29] = 1;	doodle_right_transparency_texture[75][30] = 1;	doodle_right_transparency_texture[75][31] = 1;	doodle_right_transparency_texture[75][32] = 1;	doodle_right_transparency_texture[75][33] = 1;	doodle_right_transparency_texture[75][34] = 1;	doodle_right_transparency_texture[75][35] = 1;	doodle_right_transparency_texture[75][36] = 1;	doodle_right_transparency_texture[75][37] = 1;	doodle_right_transparency_texture[75][38] = 1;	doodle_right_transparency_texture[75][39] = 1;	doodle_right_transparency_texture[75][40] = 1;	doodle_right_transparency_texture[75][41] = 1;	doodle_right_transparency_texture[75][42] = 1;	doodle_right_transparency_texture[75][43] = 1;	doodle_right_transparency_texture[75][44] = 1;	doodle_right_transparency_texture[75][45] = 1;	doodle_right_transparency_texture[75][46] = 1;	doodle_right_transparency_texture[75][47] = 1;	doodle_right_transparency_texture[75][48] = 1;	doodle_right_transparency_texture[75][49] = 1;	doodle_right_transparency_texture[75][50] = 1;	doodle_right_transparency_texture[75][51] = 1;	doodle_right_transparency_texture[75][52] = 1;	doodle_right_transparency_texture[75][53] = 1;	doodle_right_transparency_texture[75][54] = 1;	doodle_right_transparency_texture[75][55] = 1;	doodle_right_transparency_texture[75][56] = 1;	doodle_right_transparency_texture[75][57] = 1;	doodle_right_transparency_texture[75][58] = 1;	doodle_right_transparency_texture[75][59] = 1;	doodle_right_transparency_texture[75][60] = 1;	doodle_right_transparency_texture[75][61] = 1;	doodle_right_transparency_texture[75][62] = 1;	doodle_right_transparency_texture[75][63] = 1;	doodle_right_transparency_texture[75][64] = 1;	doodle_right_transparency_texture[75][65] = 1;	doodle_right_transparency_texture[75][66] = 1;	doodle_right_transparency_texture[75][67] = 1;	doodle_right_transparency_texture[75][68] = 1;	doodle_right_transparency_texture[75][69] = 1;	doodle_right_transparency_texture[75][70] = 1;	doodle_right_transparency_texture[75][71] = 1;	doodle_right_transparency_texture[75][72] = 1;	doodle_right_transparency_texture[75][73] = 1;	doodle_right_transparency_texture[75][74] = 1;	doodle_right_transparency_texture[75][75] = 1;	doodle_right_transparency_texture[75][76] = 1;	doodle_right_transparency_texture[75][77] = 1;	doodle_right_transparency_texture[75][78] = 1;	doodle_right_transparency_texture[75][79] = 1;	doodle_right_transparency_texture[76][0] = 1;	doodle_right_transparency_texture[76][1] = 1;	doodle_right_transparency_texture[76][2] = 1;	doodle_right_transparency_texture[76][3] = 1;	doodle_right_transparency_texture[76][4] = 1;	doodle_right_transparency_texture[76][5] = 1;	doodle_right_transparency_texture[76][6] = 1;	doodle_right_transparency_texture[76][7] = 1;	doodle_right_transparency_texture[76][8] = 1;	doodle_right_transparency_texture[76][9] = 1;	doodle_right_transparency_texture[76][10] = 1;	doodle_right_transparency_texture[76][11] = 1;	doodle_right_transparency_texture[76][12] = 1;	doodle_right_transparency_texture[76][13] = 1;	doodle_right_transparency_texture[76][14] = 1;	doodle_right_transparency_texture[76][15] = 1;	doodle_right_transparency_texture[76][16] = 1;	doodle_right_transparency_texture[76][17] = 1;	doodle_right_transparency_texture[76][18] = 1;	doodle_right_transparency_texture[76][19] = 1;	doodle_right_transparency_texture[76][20] = 1;	doodle_right_transparency_texture[76][21] = 1;	doodle_right_transparency_texture[76][22] = 1;	doodle_right_transparency_texture[76][23] = 1;	doodle_right_transparency_texture[76][24] = 1;	doodle_right_transparency_texture[76][25] = 1;	doodle_right_transparency_texture[76][26] = 1;	doodle_right_transparency_texture[76][27] = 1;	doodle_right_transparency_texture[76][28] = 1;	doodle_right_transparency_texture[76][29] = 1;	doodle_right_transparency_texture[76][30] = 1;	doodle_right_transparency_texture[76][31] = 1;	doodle_right_transparency_texture[76][32] = 1;	doodle_right_transparency_texture[76][33] = 1;	doodle_right_transparency_texture[76][34] = 1;	doodle_right_transparency_texture[76][35] = 1;	doodle_right_transparency_texture[76][36] = 1;	doodle_right_transparency_texture[76][37] = 1;	doodle_right_transparency_texture[76][38] = 1;	doodle_right_transparency_texture[76][39] = 1;	doodle_right_transparency_texture[76][40] = 1;	doodle_right_transparency_texture[76][41] = 1;	doodle_right_transparency_texture[76][42] = 1;	doodle_right_transparency_texture[76][43] = 1;	doodle_right_transparency_texture[76][44] = 1;	doodle_right_transparency_texture[76][45] = 1;	doodle_right_transparency_texture[76][46] = 1;	doodle_right_transparency_texture[76][47] = 1;	doodle_right_transparency_texture[76][48] = 1;	doodle_right_transparency_texture[76][49] = 1;	doodle_right_transparency_texture[76][50] = 1;	doodle_right_transparency_texture[76][51] = 1;	doodle_right_transparency_texture[76][52] = 1;	doodle_right_transparency_texture[76][53] = 1;	doodle_right_transparency_texture[76][54] = 1;	doodle_right_transparency_texture[76][55] = 1;	doodle_right_transparency_texture[76][56] = 1;	doodle_right_transparency_texture[76][57] = 1;	doodle_right_transparency_texture[76][58] = 1;	doodle_right_transparency_texture[76][59] = 1;	doodle_right_transparency_texture[76][60] = 1;	doodle_right_transparency_texture[76][61] = 1;	doodle_right_transparency_texture[76][62] = 1;	doodle_right_transparency_texture[76][63] = 1;	doodle_right_transparency_texture[76][64] = 1;	doodle_right_transparency_texture[76][65] = 1;	doodle_right_transparency_texture[76][66] = 1;	doodle_right_transparency_texture[76][67] = 1;	doodle_right_transparency_texture[76][68] = 1;	doodle_right_transparency_texture[76][69] = 1;	doodle_right_transparency_texture[76][70] = 1;	doodle_right_transparency_texture[76][71] = 1;	doodle_right_transparency_texture[76][72] = 1;	doodle_right_transparency_texture[76][73] = 1;	doodle_right_transparency_texture[76][74] = 1;	doodle_right_transparency_texture[76][75] = 1;	doodle_right_transparency_texture[76][76] = 1;	doodle_right_transparency_texture[76][77] = 1;	doodle_right_transparency_texture[76][78] = 1;	doodle_right_transparency_texture[76][79] = 1;	doodle_right_transparency_texture[77][0] = 1;	doodle_right_transparency_texture[77][1] = 1;	doodle_right_transparency_texture[77][2] = 1;	doodle_right_transparency_texture[77][3] = 1;	doodle_right_transparency_texture[77][4] = 1;	doodle_right_transparency_texture[77][5] = 1;	doodle_right_transparency_texture[77][6] = 1;	doodle_right_transparency_texture[77][7] = 1;	doodle_right_transparency_texture[77][8] = 1;	doodle_right_transparency_texture[77][9] = 1;	doodle_right_transparency_texture[77][10] = 1;	doodle_right_transparency_texture[77][11] = 1;	doodle_right_transparency_texture[77][12] = 1;	doodle_right_transparency_texture[77][13] = 1;	doodle_right_transparency_texture[77][14] = 1;	doodle_right_transparency_texture[77][15] = 1;	doodle_right_transparency_texture[77][16] = 1;	doodle_right_transparency_texture[77][17] = 1;	doodle_right_transparency_texture[77][18] = 1;	doodle_right_transparency_texture[77][19] = 1;	doodle_right_transparency_texture[77][20] = 1;	doodle_right_transparency_texture[77][21] = 1;	doodle_right_transparency_texture[77][22] = 1;	doodle_right_transparency_texture[77][23] = 1;	doodle_right_transparency_texture[77][24] = 1;	doodle_right_transparency_texture[77][25] = 1;	doodle_right_transparency_texture[77][26] = 1;	doodle_right_transparency_texture[77][27] = 1;	doodle_right_transparency_texture[77][28] = 1;	doodle_right_transparency_texture[77][29] = 1;	doodle_right_transparency_texture[77][30] = 1;	doodle_right_transparency_texture[77][31] = 1;	doodle_right_transparency_texture[77][32] = 1;	doodle_right_transparency_texture[77][33] = 1;	doodle_right_transparency_texture[77][34] = 1;	doodle_right_transparency_texture[77][35] = 1;	doodle_right_transparency_texture[77][36] = 1;	doodle_right_transparency_texture[77][37] = 1;	doodle_right_transparency_texture[77][38] = 1;	doodle_right_transparency_texture[77][39] = 1;	doodle_right_transparency_texture[77][40] = 1;	doodle_right_transparency_texture[77][41] = 1;	doodle_right_transparency_texture[77][42] = 1;	doodle_right_transparency_texture[77][43] = 1;	doodle_right_transparency_texture[77][44] = 1;	doodle_right_transparency_texture[77][45] = 1;	doodle_right_transparency_texture[77][46] = 1;	doodle_right_transparency_texture[77][47] = 1;	doodle_right_transparency_texture[77][48] = 1;	doodle_right_transparency_texture[77][49] = 1;	doodle_right_transparency_texture[77][50] = 1;	doodle_right_transparency_texture[77][51] = 1;	doodle_right_transparency_texture[77][52] = 1;	doodle_right_transparency_texture[77][53] = 1;	doodle_right_transparency_texture[77][54] = 1;	doodle_right_transparency_texture[77][55] = 1;	doodle_right_transparency_texture[77][56] = 1;	doodle_right_transparency_texture[77][57] = 1;	doodle_right_transparency_texture[77][58] = 1;	doodle_right_transparency_texture[77][59] = 1;	doodle_right_transparency_texture[77][60] = 1;	doodle_right_transparency_texture[77][61] = 1;	doodle_right_transparency_texture[77][62] = 1;	doodle_right_transparency_texture[77][63] = 1;	doodle_right_transparency_texture[77][64] = 1;	doodle_right_transparency_texture[77][65] = 1;	doodle_right_transparency_texture[77][66] = 1;	doodle_right_transparency_texture[77][67] = 1;	doodle_right_transparency_texture[77][68] = 1;	doodle_right_transparency_texture[77][69] = 1;	doodle_right_transparency_texture[77][70] = 1;	doodle_right_transparency_texture[77][71] = 1;	doodle_right_transparency_texture[77][72] = 1;	doodle_right_transparency_texture[77][73] = 1;	doodle_right_transparency_texture[77][74] = 1;	doodle_right_transparency_texture[77][75] = 1;	doodle_right_transparency_texture[77][76] = 1;	doodle_right_transparency_texture[77][77] = 1;	doodle_right_transparency_texture[77][78] = 1;	doodle_right_transparency_texture[77][79] = 1;	doodle_right_transparency_texture[78][0] = 1;	doodle_right_transparency_texture[78][1] = 1;	doodle_right_transparency_texture[78][2] = 1;	doodle_right_transparency_texture[78][3] = 1;	doodle_right_transparency_texture[78][4] = 1;	doodle_right_transparency_texture[78][5] = 1;	doodle_right_transparency_texture[78][6] = 1;	doodle_right_transparency_texture[78][7] = 1;	doodle_right_transparency_texture[78][8] = 1;	doodle_right_transparency_texture[78][9] = 1;	doodle_right_transparency_texture[78][10] = 1;	doodle_right_transparency_texture[78][11] = 1;	doodle_right_transparency_texture[78][12] = 1;	doodle_right_transparency_texture[78][13] = 1;	doodle_right_transparency_texture[78][14] = 1;	doodle_right_transparency_texture[78][15] = 1;	doodle_right_transparency_texture[78][16] = 1;	doodle_right_transparency_texture[78][17] = 1;	doodle_right_transparency_texture[78][18] = 1;	doodle_right_transparency_texture[78][19] = 1;	doodle_right_transparency_texture[78][20] = 1;	doodle_right_transparency_texture[78][21] = 1;	doodle_right_transparency_texture[78][22] = 1;	doodle_right_transparency_texture[78][23] = 1;	doodle_right_transparency_texture[78][24] = 1;	doodle_right_transparency_texture[78][25] = 1;	doodle_right_transparency_texture[78][26] = 1;	doodle_right_transparency_texture[78][27] = 1;	doodle_right_transparency_texture[78][28] = 1;	doodle_right_transparency_texture[78][29] = 1;	doodle_right_transparency_texture[78][30] = 1;	doodle_right_transparency_texture[78][31] = 1;	doodle_right_transparency_texture[78][32] = 1;	doodle_right_transparency_texture[78][33] = 1;	doodle_right_transparency_texture[78][34] = 1;	doodle_right_transparency_texture[78][35] = 1;	doodle_right_transparency_texture[78][36] = 1;	doodle_right_transparency_texture[78][37] = 1;	doodle_right_transparency_texture[78][38] = 1;	doodle_right_transparency_texture[78][39] = 1;	doodle_right_transparency_texture[78][40] = 1;	doodle_right_transparency_texture[78][41] = 1;	doodle_right_transparency_texture[78][42] = 1;	doodle_right_transparency_texture[78][43] = 1;	doodle_right_transparency_texture[78][44] = 1;	doodle_right_transparency_texture[78][45] = 1;	doodle_right_transparency_texture[78][46] = 1;	doodle_right_transparency_texture[78][47] = 1;	doodle_right_transparency_texture[78][48] = 1;	doodle_right_transparency_texture[78][49] = 1;	doodle_right_transparency_texture[78][50] = 1;	doodle_right_transparency_texture[78][51] = 1;	doodle_right_transparency_texture[78][52] = 1;	doodle_right_transparency_texture[78][53] = 1;	doodle_right_transparency_texture[78][54] = 1;	doodle_right_transparency_texture[78][55] = 1;	doodle_right_transparency_texture[78][56] = 1;	doodle_right_transparency_texture[78][57] = 1;	doodle_right_transparency_texture[78][58] = 1;	doodle_right_transparency_texture[78][59] = 1;	doodle_right_transparency_texture[78][60] = 1;	doodle_right_transparency_texture[78][61] = 1;	doodle_right_transparency_texture[78][62] = 1;	doodle_right_transparency_texture[78][63] = 1;	doodle_right_transparency_texture[78][64] = 1;	doodle_right_transparency_texture[78][65] = 1;	doodle_right_transparency_texture[78][66] = 1;	doodle_right_transparency_texture[78][67] = 1;	doodle_right_transparency_texture[78][68] = 1;	doodle_right_transparency_texture[78][69] = 1;	doodle_right_transparency_texture[78][70] = 1;	doodle_right_transparency_texture[78][71] = 1;	doodle_right_transparency_texture[78][72] = 1;	doodle_right_transparency_texture[78][73] = 1;	doodle_right_transparency_texture[78][74] = 1;	doodle_right_transparency_texture[78][75] = 1;	doodle_right_transparency_texture[78][76] = 1;	doodle_right_transparency_texture[78][77] = 1;	doodle_right_transparency_texture[78][78] = 1;	doodle_right_transparency_texture[78][79] = 1;	doodle_right_transparency_texture[79][0] = 1;	doodle_right_transparency_texture[79][1] = 1;	doodle_right_transparency_texture[79][2] = 1;	doodle_right_transparency_texture[79][3] = 1;	doodle_right_transparency_texture[79][4] = 1;	doodle_right_transparency_texture[79][5] = 1;	doodle_right_transparency_texture[79][6] = 1;	doodle_right_transparency_texture[79][7] = 1;	doodle_right_transparency_texture[79][8] = 1;	doodle_right_transparency_texture[79][9] = 1;	doodle_right_transparency_texture[79][10] = 1;	doodle_right_transparency_texture[79][11] = 1;	doodle_right_transparency_texture[79][12] = 1;	doodle_right_transparency_texture[79][13] = 1;	doodle_right_transparency_texture[79][14] = 1;	doodle_right_transparency_texture[79][15] = 1;	doodle_right_transparency_texture[79][16] = 1;	doodle_right_transparency_texture[79][17] = 1;	doodle_right_transparency_texture[79][18] = 1;	doodle_right_transparency_texture[79][19] = 1;	doodle_right_transparency_texture[79][20] = 1;	doodle_right_transparency_texture[79][21] = 1;	doodle_right_transparency_texture[79][22] = 1;	doodle_right_transparency_texture[79][23] = 1;	doodle_right_transparency_texture[79][24] = 1;	doodle_right_transparency_texture[79][25] = 1;	doodle_right_transparency_texture[79][26] = 1;	doodle_right_transparency_texture[79][27] = 1;	doodle_right_transparency_texture[79][28] = 1;	doodle_right_transparency_texture[79][29] = 1;	doodle_right_transparency_texture[79][30] = 1;	doodle_right_transparency_texture[79][31] = 1;	doodle_right_transparency_texture[79][32] = 1;	doodle_right_transparency_texture[79][33] = 1;	doodle_right_transparency_texture[79][34] = 1;	doodle_right_transparency_texture[79][35] = 1;	doodle_right_transparency_texture[79][36] = 1;	doodle_right_transparency_texture[79][37] = 1;	doodle_right_transparency_texture[79][38] = 1;	doodle_right_transparency_texture[79][39] = 1;	doodle_right_transparency_texture[79][40] = 1;	doodle_right_transparency_texture[79][41] = 1;	doodle_right_transparency_texture[79][42] = 1;	doodle_right_transparency_texture[79][43] = 1;	doodle_right_transparency_texture[79][44] = 1;	doodle_right_transparency_texture[79][45] = 1;	doodle_right_transparency_texture[79][46] = 1;	doodle_right_transparency_texture[79][47] = 1;	doodle_right_transparency_texture[79][48] = 1;	doodle_right_transparency_texture[79][49] = 1;	doodle_right_transparency_texture[79][50] = 1;	doodle_right_transparency_texture[79][51] = 1;	doodle_right_transparency_texture[79][52] = 1;	doodle_right_transparency_texture[79][53] = 1;	doodle_right_transparency_texture[79][54] = 1;	doodle_right_transparency_texture[79][55] = 1;	doodle_right_transparency_texture[79][56] = 1;	doodle_right_transparency_texture[79][57] = 1;	doodle_right_transparency_texture[79][58] = 1;	doodle_right_transparency_texture[79][59] = 1;	doodle_right_transparency_texture[79][60] = 1;	doodle_right_transparency_texture[79][61] = 1;	doodle_right_transparency_texture[79][62] = 1;	doodle_right_transparency_texture[79][63] = 1;	doodle_right_transparency_texture[79][64] = 1;	doodle_right_transparency_texture[79][65] = 1;	doodle_right_transparency_texture[79][66] = 1;	doodle_right_transparency_texture[79][67] = 1;	doodle_right_transparency_texture[79][68] = 1;	doodle_right_transparency_texture[79][69] = 1;	doodle_right_transparency_texture[79][70] = 1;	doodle_right_transparency_texture[79][71] = 1;	doodle_right_transparency_texture[79][72] = 1;	doodle_right_transparency_texture[79][73] = 1;	doodle_right_transparency_texture[79][74] = 1;	doodle_right_transparency_texture[79][75] = 1;	doodle_right_transparency_texture[79][76] = 1;	doodle_right_transparency_texture[79][77] = 1;	doodle_right_transparency_texture[79][78] = 1;	doodle_right_transparency_texture[79][79] = 1;
		doodle_left_texture[0][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[0][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[1][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[2][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[3][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[4][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[5][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[6][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[7][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[8][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[9][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[10][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[11][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[12][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[12][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[13][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[13][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[14][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[14][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[15][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[15][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[16][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[16][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[17][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[17][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[18][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[18][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[19][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[19][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[20][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[20][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[21][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[21][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[22][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[22][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[23][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[23][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[24][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[24][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[25][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[25][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[26][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[26][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[27][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[27][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][8] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][9] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][10] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][11] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][16] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][17] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][18] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][19] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][20] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][21] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][22] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][23] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][24] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][25] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][26] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][27] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[28][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[28][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][8] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][9] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][10] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][11] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][16] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][17] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][18] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][19] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][20] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][21] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][22] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][23] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][24] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][25] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][26] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][27] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[29][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[29][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][8] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][9] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][10] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][11] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][16] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][17] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][18] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][19] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][20] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][21] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][22] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][23] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][24] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][25] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][26] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][27] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[30][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[30][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][8] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][9] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][10] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][11] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][16] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][17] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][18] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][19] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][20] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][21] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][22] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][23] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][24] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][25] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][26] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][27] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[31][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[31][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[32][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[32][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[33][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[33][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[34][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[34][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][28] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][29] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][30] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][31] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[35][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[35][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[36][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[36][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[37][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[37][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[38][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[38][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[39][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[39][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[40][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[40][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[41][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[41][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[42][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[42][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[43][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[43][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[44][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[45][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[46][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[47][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[48][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[48][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[49][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[49][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[50][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[50][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[51][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[51][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[52][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[52][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[53][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[53][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[54][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[54][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][32] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][33] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][34] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][35] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][36] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][37] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][38] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][39] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][40] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][41] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][42] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][43] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][44] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][45] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][46] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][47] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][48] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][49] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][50] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][51] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][52] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][53] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][54] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][55] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][56] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][57] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][58] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][59] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][60] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][61] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][62] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][63] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][64] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][65] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][66] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][67] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][68] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][69] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][70] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][71] = {4'b0, 4'b1111, 4'b0};	doodle_left_texture[55][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[55][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[56][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[57][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[58][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[59][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[60][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[61][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[62][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[63][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[64][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[65][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[66][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[67][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[68][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[69][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[70][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[71][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[72][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[73][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[74][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[75][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[76][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[77][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[78][79] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][0] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][1] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][2] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][3] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][4] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][5] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][6] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][7] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][8] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][9] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][10] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][11] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][12] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][13] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][14] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][15] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][16] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][17] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][18] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][19] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][20] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][21] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][22] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][23] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][24] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][25] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][26] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][27] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][28] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][29] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][30] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][31] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][32] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][33] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][34] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][35] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][36] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][37] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][38] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][39] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][40] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][41] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][42] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][43] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][44] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][45] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][46] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][47] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][48] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][49] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][50] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][51] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][52] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][53] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][54] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][55] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][56] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][57] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][58] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][59] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][60] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][61] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][62] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][63] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][64] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][65] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][66] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][67] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][68] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][69] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][70] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][71] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][72] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][73] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][74] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][75] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][76] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][77] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][78] = {4'b0, 4'b0, 4'b0};	doodle_left_texture[79][79] = {4'b0, 4'b0, 4'b0};
		doodle_left_transparency_texture[0][0] = 1;	doodle_left_transparency_texture[0][1] = 1;	doodle_left_transparency_texture[0][2] = 1;	doodle_left_transparency_texture[0][3] = 1;	doodle_left_transparency_texture[0][4] = 1;	doodle_left_transparency_texture[0][5] = 1;	doodle_left_transparency_texture[0][6] = 1;	doodle_left_transparency_texture[0][7] = 1;	doodle_left_transparency_texture[0][8] = 1;	doodle_left_transparency_texture[0][9] = 1;	doodle_left_transparency_texture[0][10] = 1;	doodle_left_transparency_texture[0][11] = 1;	doodle_left_transparency_texture[0][12] = 1;	doodle_left_transparency_texture[0][13] = 1;	doodle_left_transparency_texture[0][14] = 1;	doodle_left_transparency_texture[0][15] = 1;	doodle_left_transparency_texture[0][16] = 1;	doodle_left_transparency_texture[0][17] = 1;	doodle_left_transparency_texture[0][18] = 1;	doodle_left_transparency_texture[0][19] = 1;	doodle_left_transparency_texture[0][20] = 1;	doodle_left_transparency_texture[0][21] = 1;	doodle_left_transparency_texture[0][22] = 1;	doodle_left_transparency_texture[0][23] = 1;	doodle_left_transparency_texture[0][24] = 1;	doodle_left_transparency_texture[0][25] = 1;	doodle_left_transparency_texture[0][26] = 1;	doodle_left_transparency_texture[0][27] = 1;	doodle_left_transparency_texture[0][28] = 1;	doodle_left_transparency_texture[0][29] = 1;	doodle_left_transparency_texture[0][30] = 1;	doodle_left_transparency_texture[0][31] = 1;	doodle_left_transparency_texture[0][32] = 1;	doodle_left_transparency_texture[0][33] = 1;	doodle_left_transparency_texture[0][34] = 1;	doodle_left_transparency_texture[0][35] = 1;	doodle_left_transparency_texture[0][36] = 1;	doodle_left_transparency_texture[0][37] = 1;	doodle_left_transparency_texture[0][38] = 1;	doodle_left_transparency_texture[0][39] = 1;	doodle_left_transparency_texture[0][40] = 1;	doodle_left_transparency_texture[0][41] = 1;	doodle_left_transparency_texture[0][42] = 1;	doodle_left_transparency_texture[0][43] = 1;	doodle_left_transparency_texture[0][44] = 1;	doodle_left_transparency_texture[0][45] = 1;	doodle_left_transparency_texture[0][46] = 1;	doodle_left_transparency_texture[0][47] = 1;	doodle_left_transparency_texture[0][48] = 1;	doodle_left_transparency_texture[0][49] = 1;	doodle_left_transparency_texture[0][50] = 1;	doodle_left_transparency_texture[0][51] = 1;	doodle_left_transparency_texture[0][52] = 1;	doodle_left_transparency_texture[0][53] = 1;	doodle_left_transparency_texture[0][54] = 1;	doodle_left_transparency_texture[0][55] = 1;	doodle_left_transparency_texture[0][56] = 1;	doodle_left_transparency_texture[0][57] = 1;	doodle_left_transparency_texture[0][58] = 1;	doodle_left_transparency_texture[0][59] = 1;	doodle_left_transparency_texture[0][60] = 1;	doodle_left_transparency_texture[0][61] = 1;	doodle_left_transparency_texture[0][62] = 1;	doodle_left_transparency_texture[0][63] = 1;	doodle_left_transparency_texture[0][64] = 1;	doodle_left_transparency_texture[0][65] = 1;	doodle_left_transparency_texture[0][66] = 1;	doodle_left_transparency_texture[0][67] = 1;	doodle_left_transparency_texture[0][68] = 1;	doodle_left_transparency_texture[0][69] = 1;	doodle_left_transparency_texture[0][70] = 1;	doodle_left_transparency_texture[0][71] = 1;	doodle_left_transparency_texture[0][72] = 1;	doodle_left_transparency_texture[0][73] = 1;	doodle_left_transparency_texture[0][74] = 1;	doodle_left_transparency_texture[0][75] = 1;	doodle_left_transparency_texture[0][76] = 1;	doodle_left_transparency_texture[0][77] = 1;	doodle_left_transparency_texture[0][78] = 1;	doodle_left_transparency_texture[0][79] = 1;	doodle_left_transparency_texture[1][0] = 1;	doodle_left_transparency_texture[1][1] = 1;	doodle_left_transparency_texture[1][2] = 1;	doodle_left_transparency_texture[1][3] = 1;	doodle_left_transparency_texture[1][4] = 1;	doodle_left_transparency_texture[1][5] = 1;	doodle_left_transparency_texture[1][6] = 1;	doodle_left_transparency_texture[1][7] = 1;	doodle_left_transparency_texture[1][8] = 1;	doodle_left_transparency_texture[1][9] = 1;	doodle_left_transparency_texture[1][10] = 1;	doodle_left_transparency_texture[1][11] = 1;	doodle_left_transparency_texture[1][12] = 1;	doodle_left_transparency_texture[1][13] = 1;	doodle_left_transparency_texture[1][14] = 1;	doodle_left_transparency_texture[1][15] = 1;	doodle_left_transparency_texture[1][16] = 1;	doodle_left_transparency_texture[1][17] = 1;	doodle_left_transparency_texture[1][18] = 1;	doodle_left_transparency_texture[1][19] = 1;	doodle_left_transparency_texture[1][20] = 1;	doodle_left_transparency_texture[1][21] = 1;	doodle_left_transparency_texture[1][22] = 1;	doodle_left_transparency_texture[1][23] = 1;	doodle_left_transparency_texture[1][24] = 1;	doodle_left_transparency_texture[1][25] = 1;	doodle_left_transparency_texture[1][26] = 1;	doodle_left_transparency_texture[1][27] = 1;	doodle_left_transparency_texture[1][28] = 1;	doodle_left_transparency_texture[1][29] = 1;	doodle_left_transparency_texture[1][30] = 1;	doodle_left_transparency_texture[1][31] = 1;	doodle_left_transparency_texture[1][32] = 1;	doodle_left_transparency_texture[1][33] = 1;	doodle_left_transparency_texture[1][34] = 1;	doodle_left_transparency_texture[1][35] = 1;	doodle_left_transparency_texture[1][36] = 1;	doodle_left_transparency_texture[1][37] = 1;	doodle_left_transparency_texture[1][38] = 1;	doodle_left_transparency_texture[1][39] = 1;	doodle_left_transparency_texture[1][40] = 1;	doodle_left_transparency_texture[1][41] = 1;	doodle_left_transparency_texture[1][42] = 1;	doodle_left_transparency_texture[1][43] = 1;	doodle_left_transparency_texture[1][44] = 1;	doodle_left_transparency_texture[1][45] = 1;	doodle_left_transparency_texture[1][46] = 1;	doodle_left_transparency_texture[1][47] = 1;	doodle_left_transparency_texture[1][48] = 1;	doodle_left_transparency_texture[1][49] = 1;	doodle_left_transparency_texture[1][50] = 1;	doodle_left_transparency_texture[1][51] = 1;	doodle_left_transparency_texture[1][52] = 1;	doodle_left_transparency_texture[1][53] = 1;	doodle_left_transparency_texture[1][54] = 1;	doodle_left_transparency_texture[1][55] = 1;	doodle_left_transparency_texture[1][56] = 1;	doodle_left_transparency_texture[1][57] = 1;	doodle_left_transparency_texture[1][58] = 1;	doodle_left_transparency_texture[1][59] = 1;	doodle_left_transparency_texture[1][60] = 1;	doodle_left_transparency_texture[1][61] = 1;	doodle_left_transparency_texture[1][62] = 1;	doodle_left_transparency_texture[1][63] = 1;	doodle_left_transparency_texture[1][64] = 1;	doodle_left_transparency_texture[1][65] = 1;	doodle_left_transparency_texture[1][66] = 1;	doodle_left_transparency_texture[1][67] = 1;	doodle_left_transparency_texture[1][68] = 1;	doodle_left_transparency_texture[1][69] = 1;	doodle_left_transparency_texture[1][70] = 1;	doodle_left_transparency_texture[1][71] = 1;	doodle_left_transparency_texture[1][72] = 1;	doodle_left_transparency_texture[1][73] = 1;	doodle_left_transparency_texture[1][74] = 1;	doodle_left_transparency_texture[1][75] = 1;	doodle_left_transparency_texture[1][76] = 1;	doodle_left_transparency_texture[1][77] = 1;	doodle_left_transparency_texture[1][78] = 1;	doodle_left_transparency_texture[1][79] = 1;	doodle_left_transparency_texture[2][0] = 1;	doodle_left_transparency_texture[2][1] = 1;	doodle_left_transparency_texture[2][2] = 1;	doodle_left_transparency_texture[2][3] = 1;	doodle_left_transparency_texture[2][4] = 1;	doodle_left_transparency_texture[2][5] = 1;	doodle_left_transparency_texture[2][6] = 1;	doodle_left_transparency_texture[2][7] = 1;	doodle_left_transparency_texture[2][8] = 1;	doodle_left_transparency_texture[2][9] = 1;	doodle_left_transparency_texture[2][10] = 1;	doodle_left_transparency_texture[2][11] = 1;	doodle_left_transparency_texture[2][12] = 1;	doodle_left_transparency_texture[2][13] = 1;	doodle_left_transparency_texture[2][14] = 1;	doodle_left_transparency_texture[2][15] = 1;	doodle_left_transparency_texture[2][16] = 1;	doodle_left_transparency_texture[2][17] = 1;	doodle_left_transparency_texture[2][18] = 1;	doodle_left_transparency_texture[2][19] = 1;	doodle_left_transparency_texture[2][20] = 1;	doodle_left_transparency_texture[2][21] = 1;	doodle_left_transparency_texture[2][22] = 1;	doodle_left_transparency_texture[2][23] = 1;	doodle_left_transparency_texture[2][24] = 1;	doodle_left_transparency_texture[2][25] = 1;	doodle_left_transparency_texture[2][26] = 1;	doodle_left_transparency_texture[2][27] = 1;	doodle_left_transparency_texture[2][28] = 1;	doodle_left_transparency_texture[2][29] = 1;	doodle_left_transparency_texture[2][30] = 1;	doodle_left_transparency_texture[2][31] = 1;	doodle_left_transparency_texture[2][32] = 1;	doodle_left_transparency_texture[2][33] = 1;	doodle_left_transparency_texture[2][34] = 1;	doodle_left_transparency_texture[2][35] = 1;	doodle_left_transparency_texture[2][36] = 1;	doodle_left_transparency_texture[2][37] = 1;	doodle_left_transparency_texture[2][38] = 1;	doodle_left_transparency_texture[2][39] = 1;	doodle_left_transparency_texture[2][40] = 1;	doodle_left_transparency_texture[2][41] = 1;	doodle_left_transparency_texture[2][42] = 1;	doodle_left_transparency_texture[2][43] = 1;	doodle_left_transparency_texture[2][44] = 1;	doodle_left_transparency_texture[2][45] = 1;	doodle_left_transparency_texture[2][46] = 1;	doodle_left_transparency_texture[2][47] = 1;	doodle_left_transparency_texture[2][48] = 1;	doodle_left_transparency_texture[2][49] = 1;	doodle_left_transparency_texture[2][50] = 1;	doodle_left_transparency_texture[2][51] = 1;	doodle_left_transparency_texture[2][52] = 1;	doodle_left_transparency_texture[2][53] = 1;	doodle_left_transparency_texture[2][54] = 1;	doodle_left_transparency_texture[2][55] = 1;	doodle_left_transparency_texture[2][56] = 1;	doodle_left_transparency_texture[2][57] = 1;	doodle_left_transparency_texture[2][58] = 1;	doodle_left_transparency_texture[2][59] = 1;	doodle_left_transparency_texture[2][60] = 1;	doodle_left_transparency_texture[2][61] = 1;	doodle_left_transparency_texture[2][62] = 1;	doodle_left_transparency_texture[2][63] = 1;	doodle_left_transparency_texture[2][64] = 1;	doodle_left_transparency_texture[2][65] = 1;	doodle_left_transparency_texture[2][66] = 1;	doodle_left_transparency_texture[2][67] = 1;	doodle_left_transparency_texture[2][68] = 1;	doodle_left_transparency_texture[2][69] = 1;	doodle_left_transparency_texture[2][70] = 1;	doodle_left_transparency_texture[2][71] = 1;	doodle_left_transparency_texture[2][72] = 1;	doodle_left_transparency_texture[2][73] = 1;	doodle_left_transparency_texture[2][74] = 1;	doodle_left_transparency_texture[2][75] = 1;	doodle_left_transparency_texture[2][76] = 1;	doodle_left_transparency_texture[2][77] = 1;	doodle_left_transparency_texture[2][78] = 1;	doodle_left_transparency_texture[2][79] = 1;	doodle_left_transparency_texture[3][0] = 1;	doodle_left_transparency_texture[3][1] = 1;	doodle_left_transparency_texture[3][2] = 1;	doodle_left_transparency_texture[3][3] = 1;	doodle_left_transparency_texture[3][4] = 1;	doodle_left_transparency_texture[3][5] = 1;	doodle_left_transparency_texture[3][6] = 1;	doodle_left_transparency_texture[3][7] = 1;	doodle_left_transparency_texture[3][8] = 1;	doodle_left_transparency_texture[3][9] = 1;	doodle_left_transparency_texture[3][10] = 1;	doodle_left_transparency_texture[3][11] = 1;	doodle_left_transparency_texture[3][12] = 1;	doodle_left_transparency_texture[3][13] = 1;	doodle_left_transparency_texture[3][14] = 1;	doodle_left_transparency_texture[3][15] = 1;	doodle_left_transparency_texture[3][16] = 1;	doodle_left_transparency_texture[3][17] = 1;	doodle_left_transparency_texture[3][18] = 1;	doodle_left_transparency_texture[3][19] = 1;	doodle_left_transparency_texture[3][20] = 1;	doodle_left_transparency_texture[3][21] = 1;	doodle_left_transparency_texture[3][22] = 1;	doodle_left_transparency_texture[3][23] = 1;	doodle_left_transparency_texture[3][24] = 1;	doodle_left_transparency_texture[3][25] = 1;	doodle_left_transparency_texture[3][26] = 1;	doodle_left_transparency_texture[3][27] = 1;	doodle_left_transparency_texture[3][28] = 1;	doodle_left_transparency_texture[3][29] = 1;	doodle_left_transparency_texture[3][30] = 1;	doodle_left_transparency_texture[3][31] = 1;	doodle_left_transparency_texture[3][32] = 1;	doodle_left_transparency_texture[3][33] = 1;	doodle_left_transparency_texture[3][34] = 1;	doodle_left_transparency_texture[3][35] = 1;	doodle_left_transparency_texture[3][36] = 1;	doodle_left_transparency_texture[3][37] = 1;	doodle_left_transparency_texture[3][38] = 1;	doodle_left_transparency_texture[3][39] = 1;	doodle_left_transparency_texture[3][40] = 1;	doodle_left_transparency_texture[3][41] = 1;	doodle_left_transparency_texture[3][42] = 1;	doodle_left_transparency_texture[3][43] = 1;	doodle_left_transparency_texture[3][44] = 1;	doodle_left_transparency_texture[3][45] = 1;	doodle_left_transparency_texture[3][46] = 1;	doodle_left_transparency_texture[3][47] = 1;	doodle_left_transparency_texture[3][48] = 1;	doodle_left_transparency_texture[3][49] = 1;	doodle_left_transparency_texture[3][50] = 1;	doodle_left_transparency_texture[3][51] = 1;	doodle_left_transparency_texture[3][52] = 1;	doodle_left_transparency_texture[3][53] = 1;	doodle_left_transparency_texture[3][54] = 1;	doodle_left_transparency_texture[3][55] = 1;	doodle_left_transparency_texture[3][56] = 1;	doodle_left_transparency_texture[3][57] = 1;	doodle_left_transparency_texture[3][58] = 1;	doodle_left_transparency_texture[3][59] = 1;	doodle_left_transparency_texture[3][60] = 1;	doodle_left_transparency_texture[3][61] = 1;	doodle_left_transparency_texture[3][62] = 1;	doodle_left_transparency_texture[3][63] = 1;	doodle_left_transparency_texture[3][64] = 1;	doodle_left_transparency_texture[3][65] = 1;	doodle_left_transparency_texture[3][66] = 1;	doodle_left_transparency_texture[3][67] = 1;	doodle_left_transparency_texture[3][68] = 1;	doodle_left_transparency_texture[3][69] = 1;	doodle_left_transparency_texture[3][70] = 1;	doodle_left_transparency_texture[3][71] = 1;	doodle_left_transparency_texture[3][72] = 1;	doodle_left_transparency_texture[3][73] = 1;	doodle_left_transparency_texture[3][74] = 1;	doodle_left_transparency_texture[3][75] = 1;	doodle_left_transparency_texture[3][76] = 1;	doodle_left_transparency_texture[3][77] = 1;	doodle_left_transparency_texture[3][78] = 1;	doodle_left_transparency_texture[3][79] = 1;	doodle_left_transparency_texture[4][0] = 1;	doodle_left_transparency_texture[4][1] = 1;	doodle_left_transparency_texture[4][2] = 1;	doodle_left_transparency_texture[4][3] = 1;	doodle_left_transparency_texture[4][4] = 1;	doodle_left_transparency_texture[4][5] = 1;	doodle_left_transparency_texture[4][6] = 1;	doodle_left_transparency_texture[4][7] = 1;	doodle_left_transparency_texture[4][8] = 1;	doodle_left_transparency_texture[4][9] = 1;	doodle_left_transparency_texture[4][10] = 1;	doodle_left_transparency_texture[4][11] = 1;	doodle_left_transparency_texture[4][12] = 1;	doodle_left_transparency_texture[4][13] = 1;	doodle_left_transparency_texture[4][14] = 1;	doodle_left_transparency_texture[4][15] = 1;	doodle_left_transparency_texture[4][16] = 1;	doodle_left_transparency_texture[4][17] = 1;	doodle_left_transparency_texture[4][18] = 1;	doodle_left_transparency_texture[4][19] = 1;	doodle_left_transparency_texture[4][20] = 1;	doodle_left_transparency_texture[4][21] = 1;	doodle_left_transparency_texture[4][22] = 1;	doodle_left_transparency_texture[4][23] = 1;	doodle_left_transparency_texture[4][24] = 1;	doodle_left_transparency_texture[4][25] = 1;	doodle_left_transparency_texture[4][26] = 1;	doodle_left_transparency_texture[4][27] = 1;	doodle_left_transparency_texture[4][28] = 1;	doodle_left_transparency_texture[4][29] = 1;	doodle_left_transparency_texture[4][30] = 1;	doodle_left_transparency_texture[4][31] = 1;	doodle_left_transparency_texture[4][32] = 1;	doodle_left_transparency_texture[4][33] = 1;	doodle_left_transparency_texture[4][34] = 1;	doodle_left_transparency_texture[4][35] = 1;	doodle_left_transparency_texture[4][36] = 1;	doodle_left_transparency_texture[4][37] = 1;	doodle_left_transparency_texture[4][38] = 1;	doodle_left_transparency_texture[4][39] = 1;	doodle_left_transparency_texture[4][40] = 1;	doodle_left_transparency_texture[4][41] = 1;	doodle_left_transparency_texture[4][42] = 1;	doodle_left_transparency_texture[4][43] = 1;	doodle_left_transparency_texture[4][44] = 1;	doodle_left_transparency_texture[4][45] = 1;	doodle_left_transparency_texture[4][46] = 1;	doodle_left_transparency_texture[4][47] = 1;	doodle_left_transparency_texture[4][48] = 1;	doodle_left_transparency_texture[4][49] = 1;	doodle_left_transparency_texture[4][50] = 1;	doodle_left_transparency_texture[4][51] = 1;	doodle_left_transparency_texture[4][52] = 1;	doodle_left_transparency_texture[4][53] = 1;	doodle_left_transparency_texture[4][54] = 1;	doodle_left_transparency_texture[4][55] = 1;	doodle_left_transparency_texture[4][56] = 1;	doodle_left_transparency_texture[4][57] = 1;	doodle_left_transparency_texture[4][58] = 1;	doodle_left_transparency_texture[4][59] = 1;	doodle_left_transparency_texture[4][60] = 1;	doodle_left_transparency_texture[4][61] = 1;	doodle_left_transparency_texture[4][62] = 1;	doodle_left_transparency_texture[4][63] = 1;	doodle_left_transparency_texture[4][64] = 1;	doodle_left_transparency_texture[4][65] = 1;	doodle_left_transparency_texture[4][66] = 1;	doodle_left_transparency_texture[4][67] = 1;	doodle_left_transparency_texture[4][68] = 1;	doodle_left_transparency_texture[4][69] = 1;	doodle_left_transparency_texture[4][70] = 1;	doodle_left_transparency_texture[4][71] = 1;	doodle_left_transparency_texture[4][72] = 1;	doodle_left_transparency_texture[4][73] = 1;	doodle_left_transparency_texture[4][74] = 1;	doodle_left_transparency_texture[4][75] = 1;	doodle_left_transparency_texture[4][76] = 1;	doodle_left_transparency_texture[4][77] = 1;	doodle_left_transparency_texture[4][78] = 1;	doodle_left_transparency_texture[4][79] = 1;	doodle_left_transparency_texture[5][0] = 1;	doodle_left_transparency_texture[5][1] = 1;	doodle_left_transparency_texture[5][2] = 1;	doodle_left_transparency_texture[5][3] = 1;	doodle_left_transparency_texture[5][4] = 1;	doodle_left_transparency_texture[5][5] = 1;	doodle_left_transparency_texture[5][6] = 1;	doodle_left_transparency_texture[5][7] = 1;	doodle_left_transparency_texture[5][8] = 1;	doodle_left_transparency_texture[5][9] = 1;	doodle_left_transparency_texture[5][10] = 1;	doodle_left_transparency_texture[5][11] = 1;	doodle_left_transparency_texture[5][12] = 1;	doodle_left_transparency_texture[5][13] = 1;	doodle_left_transparency_texture[5][14] = 1;	doodle_left_transparency_texture[5][15] = 1;	doodle_left_transparency_texture[5][16] = 1;	doodle_left_transparency_texture[5][17] = 1;	doodle_left_transparency_texture[5][18] = 1;	doodle_left_transparency_texture[5][19] = 1;	doodle_left_transparency_texture[5][20] = 1;	doodle_left_transparency_texture[5][21] = 1;	doodle_left_transparency_texture[5][22] = 1;	doodle_left_transparency_texture[5][23] = 1;	doodle_left_transparency_texture[5][24] = 1;	doodle_left_transparency_texture[5][25] = 1;	doodle_left_transparency_texture[5][26] = 1;	doodle_left_transparency_texture[5][27] = 1;	doodle_left_transparency_texture[5][28] = 1;	doodle_left_transparency_texture[5][29] = 1;	doodle_left_transparency_texture[5][30] = 1;	doodle_left_transparency_texture[5][31] = 1;	doodle_left_transparency_texture[5][32] = 1;	doodle_left_transparency_texture[5][33] = 1;	doodle_left_transparency_texture[5][34] = 1;	doodle_left_transparency_texture[5][35] = 1;	doodle_left_transparency_texture[5][36] = 1;	doodle_left_transparency_texture[5][37] = 1;	doodle_left_transparency_texture[5][38] = 1;	doodle_left_transparency_texture[5][39] = 1;	doodle_left_transparency_texture[5][40] = 1;	doodle_left_transparency_texture[5][41] = 1;	doodle_left_transparency_texture[5][42] = 1;	doodle_left_transparency_texture[5][43] = 1;	doodle_left_transparency_texture[5][44] = 1;	doodle_left_transparency_texture[5][45] = 1;	doodle_left_transparency_texture[5][46] = 1;	doodle_left_transparency_texture[5][47] = 1;	doodle_left_transparency_texture[5][48] = 1;	doodle_left_transparency_texture[5][49] = 1;	doodle_left_transparency_texture[5][50] = 1;	doodle_left_transparency_texture[5][51] = 1;	doodle_left_transparency_texture[5][52] = 1;	doodle_left_transparency_texture[5][53] = 1;	doodle_left_transparency_texture[5][54] = 1;	doodle_left_transparency_texture[5][55] = 1;	doodle_left_transparency_texture[5][56] = 1;	doodle_left_transparency_texture[5][57] = 1;	doodle_left_transparency_texture[5][58] = 1;	doodle_left_transparency_texture[5][59] = 1;	doodle_left_transparency_texture[5][60] = 1;	doodle_left_transparency_texture[5][61] = 1;	doodle_left_transparency_texture[5][62] = 1;	doodle_left_transparency_texture[5][63] = 1;	doodle_left_transparency_texture[5][64] = 1;	doodle_left_transparency_texture[5][65] = 1;	doodle_left_transparency_texture[5][66] = 1;	doodle_left_transparency_texture[5][67] = 1;	doodle_left_transparency_texture[5][68] = 1;	doodle_left_transparency_texture[5][69] = 1;	doodle_left_transparency_texture[5][70] = 1;	doodle_left_transparency_texture[5][71] = 1;	doodle_left_transparency_texture[5][72] = 1;	doodle_left_transparency_texture[5][73] = 1;	doodle_left_transparency_texture[5][74] = 1;	doodle_left_transparency_texture[5][75] = 1;	doodle_left_transparency_texture[5][76] = 1;	doodle_left_transparency_texture[5][77] = 1;	doodle_left_transparency_texture[5][78] = 1;	doodle_left_transparency_texture[5][79] = 1;	doodle_left_transparency_texture[6][0] = 1;	doodle_left_transparency_texture[6][1] = 1;	doodle_left_transparency_texture[6][2] = 1;	doodle_left_transparency_texture[6][3] = 1;	doodle_left_transparency_texture[6][4] = 1;	doodle_left_transparency_texture[6][5] = 1;	doodle_left_transparency_texture[6][6] = 1;	doodle_left_transparency_texture[6][7] = 1;	doodle_left_transparency_texture[6][8] = 1;	doodle_left_transparency_texture[6][9] = 1;	doodle_left_transparency_texture[6][10] = 1;	doodle_left_transparency_texture[6][11] = 1;	doodle_left_transparency_texture[6][12] = 1;	doodle_left_transparency_texture[6][13] = 1;	doodle_left_transparency_texture[6][14] = 1;	doodle_left_transparency_texture[6][15] = 1;	doodle_left_transparency_texture[6][16] = 1;	doodle_left_transparency_texture[6][17] = 1;	doodle_left_transparency_texture[6][18] = 1;	doodle_left_transparency_texture[6][19] = 1;	doodle_left_transparency_texture[6][20] = 1;	doodle_left_transparency_texture[6][21] = 1;	doodle_left_transparency_texture[6][22] = 1;	doodle_left_transparency_texture[6][23] = 1;	doodle_left_transparency_texture[6][24] = 1;	doodle_left_transparency_texture[6][25] = 1;	doodle_left_transparency_texture[6][26] = 1;	doodle_left_transparency_texture[6][27] = 1;	doodle_left_transparency_texture[6][28] = 1;	doodle_left_transparency_texture[6][29] = 1;	doodle_left_transparency_texture[6][30] = 1;	doodle_left_transparency_texture[6][31] = 1;	doodle_left_transparency_texture[6][32] = 1;	doodle_left_transparency_texture[6][33] = 1;	doodle_left_transparency_texture[6][34] = 1;	doodle_left_transparency_texture[6][35] = 1;	doodle_left_transparency_texture[6][36] = 1;	doodle_left_transparency_texture[6][37] = 1;	doodle_left_transparency_texture[6][38] = 1;	doodle_left_transparency_texture[6][39] = 1;	doodle_left_transparency_texture[6][40] = 1;	doodle_left_transparency_texture[6][41] = 1;	doodle_left_transparency_texture[6][42] = 1;	doodle_left_transparency_texture[6][43] = 1;	doodle_left_transparency_texture[6][44] = 1;	doodle_left_transparency_texture[6][45] = 1;	doodle_left_transparency_texture[6][46] = 1;	doodle_left_transparency_texture[6][47] = 1;	doodle_left_transparency_texture[6][48] = 1;	doodle_left_transparency_texture[6][49] = 1;	doodle_left_transparency_texture[6][50] = 1;	doodle_left_transparency_texture[6][51] = 1;	doodle_left_transparency_texture[6][52] = 1;	doodle_left_transparency_texture[6][53] = 1;	doodle_left_transparency_texture[6][54] = 1;	doodle_left_transparency_texture[6][55] = 1;	doodle_left_transparency_texture[6][56] = 1;	doodle_left_transparency_texture[6][57] = 1;	doodle_left_transparency_texture[6][58] = 1;	doodle_left_transparency_texture[6][59] = 1;	doodle_left_transparency_texture[6][60] = 1;	doodle_left_transparency_texture[6][61] = 1;	doodle_left_transparency_texture[6][62] = 1;	doodle_left_transparency_texture[6][63] = 1;	doodle_left_transparency_texture[6][64] = 1;	doodle_left_transparency_texture[6][65] = 1;	doodle_left_transparency_texture[6][66] = 1;	doodle_left_transparency_texture[6][67] = 1;	doodle_left_transparency_texture[6][68] = 1;	doodle_left_transparency_texture[6][69] = 1;	doodle_left_transparency_texture[6][70] = 1;	doodle_left_transparency_texture[6][71] = 1;	doodle_left_transparency_texture[6][72] = 1;	doodle_left_transparency_texture[6][73] = 1;	doodle_left_transparency_texture[6][74] = 1;	doodle_left_transparency_texture[6][75] = 1;	doodle_left_transparency_texture[6][76] = 1;	doodle_left_transparency_texture[6][77] = 1;	doodle_left_transparency_texture[6][78] = 1;	doodle_left_transparency_texture[6][79] = 1;	doodle_left_transparency_texture[7][0] = 1;	doodle_left_transparency_texture[7][1] = 1;	doodle_left_transparency_texture[7][2] = 1;	doodle_left_transparency_texture[7][3] = 1;	doodle_left_transparency_texture[7][4] = 1;	doodle_left_transparency_texture[7][5] = 1;	doodle_left_transparency_texture[7][6] = 1;	doodle_left_transparency_texture[7][7] = 1;	doodle_left_transparency_texture[7][8] = 1;	doodle_left_transparency_texture[7][9] = 1;	doodle_left_transparency_texture[7][10] = 1;	doodle_left_transparency_texture[7][11] = 1;	doodle_left_transparency_texture[7][12] = 1;	doodle_left_transparency_texture[7][13] = 1;	doodle_left_transparency_texture[7][14] = 1;	doodle_left_transparency_texture[7][15] = 1;	doodle_left_transparency_texture[7][16] = 1;	doodle_left_transparency_texture[7][17] = 1;	doodle_left_transparency_texture[7][18] = 1;	doodle_left_transparency_texture[7][19] = 1;	doodle_left_transparency_texture[7][20] = 1;	doodle_left_transparency_texture[7][21] = 1;	doodle_left_transparency_texture[7][22] = 1;	doodle_left_transparency_texture[7][23] = 1;	doodle_left_transparency_texture[7][24] = 1;	doodle_left_transparency_texture[7][25] = 1;	doodle_left_transparency_texture[7][26] = 1;	doodle_left_transparency_texture[7][27] = 1;	doodle_left_transparency_texture[7][28] = 1;	doodle_left_transparency_texture[7][29] = 1;	doodle_left_transparency_texture[7][30] = 1;	doodle_left_transparency_texture[7][31] = 1;	doodle_left_transparency_texture[7][32] = 1;	doodle_left_transparency_texture[7][33] = 1;	doodle_left_transparency_texture[7][34] = 1;	doodle_left_transparency_texture[7][35] = 1;	doodle_left_transparency_texture[7][36] = 1;	doodle_left_transparency_texture[7][37] = 1;	doodle_left_transparency_texture[7][38] = 1;	doodle_left_transparency_texture[7][39] = 1;	doodle_left_transparency_texture[7][40] = 1;	doodle_left_transparency_texture[7][41] = 1;	doodle_left_transparency_texture[7][42] = 1;	doodle_left_transparency_texture[7][43] = 1;	doodle_left_transparency_texture[7][44] = 1;	doodle_left_transparency_texture[7][45] = 1;	doodle_left_transparency_texture[7][46] = 1;	doodle_left_transparency_texture[7][47] = 1;	doodle_left_transparency_texture[7][48] = 1;	doodle_left_transparency_texture[7][49] = 1;	doodle_left_transparency_texture[7][50] = 1;	doodle_left_transparency_texture[7][51] = 1;	doodle_left_transparency_texture[7][52] = 1;	doodle_left_transparency_texture[7][53] = 1;	doodle_left_transparency_texture[7][54] = 1;	doodle_left_transparency_texture[7][55] = 1;	doodle_left_transparency_texture[7][56] = 1;	doodle_left_transparency_texture[7][57] = 1;	doodle_left_transparency_texture[7][58] = 1;	doodle_left_transparency_texture[7][59] = 1;	doodle_left_transparency_texture[7][60] = 1;	doodle_left_transparency_texture[7][61] = 1;	doodle_left_transparency_texture[7][62] = 1;	doodle_left_transparency_texture[7][63] = 1;	doodle_left_transparency_texture[7][64] = 1;	doodle_left_transparency_texture[7][65] = 1;	doodle_left_transparency_texture[7][66] = 1;	doodle_left_transparency_texture[7][67] = 1;	doodle_left_transparency_texture[7][68] = 1;	doodle_left_transparency_texture[7][69] = 1;	doodle_left_transparency_texture[7][70] = 1;	doodle_left_transparency_texture[7][71] = 1;	doodle_left_transparency_texture[7][72] = 1;	doodle_left_transparency_texture[7][73] = 1;	doodle_left_transparency_texture[7][74] = 1;	doodle_left_transparency_texture[7][75] = 1;	doodle_left_transparency_texture[7][76] = 1;	doodle_left_transparency_texture[7][77] = 1;	doodle_left_transparency_texture[7][78] = 1;	doodle_left_transparency_texture[7][79] = 1;	doodle_left_transparency_texture[8][0] = 1;	doodle_left_transparency_texture[8][1] = 1;	doodle_left_transparency_texture[8][2] = 1;	doodle_left_transparency_texture[8][3] = 1;	doodle_left_transparency_texture[8][4] = 1;	doodle_left_transparency_texture[8][5] = 1;	doodle_left_transparency_texture[8][6] = 1;	doodle_left_transparency_texture[8][7] = 1;	doodle_left_transparency_texture[8][8] = 1;	doodle_left_transparency_texture[8][9] = 1;	doodle_left_transparency_texture[8][10] = 1;	doodle_left_transparency_texture[8][11] = 1;	doodle_left_transparency_texture[8][12] = 1;	doodle_left_transparency_texture[8][13] = 1;	doodle_left_transparency_texture[8][14] = 1;	doodle_left_transparency_texture[8][15] = 1;	doodle_left_transparency_texture[8][16] = 1;	doodle_left_transparency_texture[8][17] = 1;	doodle_left_transparency_texture[8][18] = 1;	doodle_left_transparency_texture[8][19] = 1;	doodle_left_transparency_texture[8][20] = 1;	doodle_left_transparency_texture[8][21] = 1;	doodle_left_transparency_texture[8][22] = 1;	doodle_left_transparency_texture[8][23] = 1;	doodle_left_transparency_texture[8][24] = 1;	doodle_left_transparency_texture[8][25] = 1;	doodle_left_transparency_texture[8][26] = 1;	doodle_left_transparency_texture[8][27] = 1;	doodle_left_transparency_texture[8][28] = 1;	doodle_left_transparency_texture[8][29] = 1;	doodle_left_transparency_texture[8][30] = 1;	doodle_left_transparency_texture[8][31] = 1;	doodle_left_transparency_texture[8][32] = 1;	doodle_left_transparency_texture[8][33] = 1;	doodle_left_transparency_texture[8][34] = 1;	doodle_left_transparency_texture[8][35] = 1;	doodle_left_transparency_texture[8][36] = 0;	doodle_left_transparency_texture[8][37] = 0;	doodle_left_transparency_texture[8][38] = 0;	doodle_left_transparency_texture[8][39] = 0;	doodle_left_transparency_texture[8][40] = 0;	doodle_left_transparency_texture[8][41] = 0;	doodle_left_transparency_texture[8][42] = 0;	doodle_left_transparency_texture[8][43] = 0;	doodle_left_transparency_texture[8][44] = 0;	doodle_left_transparency_texture[8][45] = 0;	doodle_left_transparency_texture[8][46] = 0;	doodle_left_transparency_texture[8][47] = 0;	doodle_left_transparency_texture[8][48] = 0;	doodle_left_transparency_texture[8][49] = 0;	doodle_left_transparency_texture[8][50] = 0;	doodle_left_transparency_texture[8][51] = 0;	doodle_left_transparency_texture[8][52] = 0;	doodle_left_transparency_texture[8][53] = 0;	doodle_left_transparency_texture[8][54] = 0;	doodle_left_transparency_texture[8][55] = 0;	doodle_left_transparency_texture[8][56] = 0;	doodle_left_transparency_texture[8][57] = 0;	doodle_left_transparency_texture[8][58] = 0;	doodle_left_transparency_texture[8][59] = 0;	doodle_left_transparency_texture[8][60] = 0;	doodle_left_transparency_texture[8][61] = 0;	doodle_left_transparency_texture[8][62] = 0;	doodle_left_transparency_texture[8][63] = 0;	doodle_left_transparency_texture[8][64] = 0;	doodle_left_transparency_texture[8][65] = 0;	doodle_left_transparency_texture[8][66] = 0;	doodle_left_transparency_texture[8][67] = 0;	doodle_left_transparency_texture[8][68] = 1;	doodle_left_transparency_texture[8][69] = 1;	doodle_left_transparency_texture[8][70] = 1;	doodle_left_transparency_texture[8][71] = 1;	doodle_left_transparency_texture[8][72] = 1;	doodle_left_transparency_texture[8][73] = 1;	doodle_left_transparency_texture[8][74] = 1;	doodle_left_transparency_texture[8][75] = 1;	doodle_left_transparency_texture[8][76] = 1;	doodle_left_transparency_texture[8][77] = 1;	doodle_left_transparency_texture[8][78] = 1;	doodle_left_transparency_texture[8][79] = 1;	doodle_left_transparency_texture[9][0] = 1;	doodle_left_transparency_texture[9][1] = 1;	doodle_left_transparency_texture[9][2] = 1;	doodle_left_transparency_texture[9][3] = 1;	doodle_left_transparency_texture[9][4] = 1;	doodle_left_transparency_texture[9][5] = 1;	doodle_left_transparency_texture[9][6] = 1;	doodle_left_transparency_texture[9][7] = 1;	doodle_left_transparency_texture[9][8] = 1;	doodle_left_transparency_texture[9][9] = 1;	doodle_left_transparency_texture[9][10] = 1;	doodle_left_transparency_texture[9][11] = 1;	doodle_left_transparency_texture[9][12] = 1;	doodle_left_transparency_texture[9][13] = 1;	doodle_left_transparency_texture[9][14] = 1;	doodle_left_transparency_texture[9][15] = 1;	doodle_left_transparency_texture[9][16] = 1;	doodle_left_transparency_texture[9][17] = 1;	doodle_left_transparency_texture[9][18] = 1;	doodle_left_transparency_texture[9][19] = 1;	doodle_left_transparency_texture[9][20] = 1;	doodle_left_transparency_texture[9][21] = 1;	doodle_left_transparency_texture[9][22] = 1;	doodle_left_transparency_texture[9][23] = 1;	doodle_left_transparency_texture[9][24] = 1;	doodle_left_transparency_texture[9][25] = 1;	doodle_left_transparency_texture[9][26] = 1;	doodle_left_transparency_texture[9][27] = 1;	doodle_left_transparency_texture[9][28] = 1;	doodle_left_transparency_texture[9][29] = 1;	doodle_left_transparency_texture[9][30] = 1;	doodle_left_transparency_texture[9][31] = 1;	doodle_left_transparency_texture[9][32] = 1;	doodle_left_transparency_texture[9][33] = 1;	doodle_left_transparency_texture[9][34] = 1;	doodle_left_transparency_texture[9][35] = 1;	doodle_left_transparency_texture[9][36] = 0;	doodle_left_transparency_texture[9][37] = 0;	doodle_left_transparency_texture[9][38] = 0;	doodle_left_transparency_texture[9][39] = 0;	doodle_left_transparency_texture[9][40] = 0;	doodle_left_transparency_texture[9][41] = 0;	doodle_left_transparency_texture[9][42] = 0;	doodle_left_transparency_texture[9][43] = 0;	doodle_left_transparency_texture[9][44] = 0;	doodle_left_transparency_texture[9][45] = 0;	doodle_left_transparency_texture[9][46] = 0;	doodle_left_transparency_texture[9][47] = 0;	doodle_left_transparency_texture[9][48] = 0;	doodle_left_transparency_texture[9][49] = 0;	doodle_left_transparency_texture[9][50] = 0;	doodle_left_transparency_texture[9][51] = 0;	doodle_left_transparency_texture[9][52] = 0;	doodle_left_transparency_texture[9][53] = 0;	doodle_left_transparency_texture[9][54] = 0;	doodle_left_transparency_texture[9][55] = 0;	doodle_left_transparency_texture[9][56] = 0;	doodle_left_transparency_texture[9][57] = 0;	doodle_left_transparency_texture[9][58] = 0;	doodle_left_transparency_texture[9][59] = 0;	doodle_left_transparency_texture[9][60] = 0;	doodle_left_transparency_texture[9][61] = 0;	doodle_left_transparency_texture[9][62] = 0;	doodle_left_transparency_texture[9][63] = 0;	doodle_left_transparency_texture[9][64] = 0;	doodle_left_transparency_texture[9][65] = 0;	doodle_left_transparency_texture[9][66] = 0;	doodle_left_transparency_texture[9][67] = 0;	doodle_left_transparency_texture[9][68] = 1;	doodle_left_transparency_texture[9][69] = 1;	doodle_left_transparency_texture[9][70] = 1;	doodle_left_transparency_texture[9][71] = 1;	doodle_left_transparency_texture[9][72] = 1;	doodle_left_transparency_texture[9][73] = 1;	doodle_left_transparency_texture[9][74] = 1;	doodle_left_transparency_texture[9][75] = 1;	doodle_left_transparency_texture[9][76] = 1;	doodle_left_transparency_texture[9][77] = 1;	doodle_left_transparency_texture[9][78] = 1;	doodle_left_transparency_texture[9][79] = 1;	doodle_left_transparency_texture[10][0] = 1;	doodle_left_transparency_texture[10][1] = 1;	doodle_left_transparency_texture[10][2] = 1;	doodle_left_transparency_texture[10][3] = 1;	doodle_left_transparency_texture[10][4] = 1;	doodle_left_transparency_texture[10][5] = 1;	doodle_left_transparency_texture[10][6] = 1;	doodle_left_transparency_texture[10][7] = 1;	doodle_left_transparency_texture[10][8] = 1;	doodle_left_transparency_texture[10][9] = 1;	doodle_left_transparency_texture[10][10] = 1;	doodle_left_transparency_texture[10][11] = 1;	doodle_left_transparency_texture[10][12] = 1;	doodle_left_transparency_texture[10][13] = 1;	doodle_left_transparency_texture[10][14] = 1;	doodle_left_transparency_texture[10][15] = 1;	doodle_left_transparency_texture[10][16] = 1;	doodle_left_transparency_texture[10][17] = 1;	doodle_left_transparency_texture[10][18] = 1;	doodle_left_transparency_texture[10][19] = 1;	doodle_left_transparency_texture[10][20] = 1;	doodle_left_transparency_texture[10][21] = 1;	doodle_left_transparency_texture[10][22] = 1;	doodle_left_transparency_texture[10][23] = 1;	doodle_left_transparency_texture[10][24] = 1;	doodle_left_transparency_texture[10][25] = 1;	doodle_left_transparency_texture[10][26] = 1;	doodle_left_transparency_texture[10][27] = 1;	doodle_left_transparency_texture[10][28] = 1;	doodle_left_transparency_texture[10][29] = 1;	doodle_left_transparency_texture[10][30] = 1;	doodle_left_transparency_texture[10][31] = 1;	doodle_left_transparency_texture[10][32] = 1;	doodle_left_transparency_texture[10][33] = 1;	doodle_left_transparency_texture[10][34] = 1;	doodle_left_transparency_texture[10][35] = 1;	doodle_left_transparency_texture[10][36] = 0;	doodle_left_transparency_texture[10][37] = 0;	doodle_left_transparency_texture[10][38] = 0;	doodle_left_transparency_texture[10][39] = 0;	doodle_left_transparency_texture[10][40] = 0;	doodle_left_transparency_texture[10][41] = 0;	doodle_left_transparency_texture[10][42] = 0;	doodle_left_transparency_texture[10][43] = 0;	doodle_left_transparency_texture[10][44] = 0;	doodle_left_transparency_texture[10][45] = 0;	doodle_left_transparency_texture[10][46] = 0;	doodle_left_transparency_texture[10][47] = 0;	doodle_left_transparency_texture[10][48] = 0;	doodle_left_transparency_texture[10][49] = 0;	doodle_left_transparency_texture[10][50] = 0;	doodle_left_transparency_texture[10][51] = 0;	doodle_left_transparency_texture[10][52] = 0;	doodle_left_transparency_texture[10][53] = 0;	doodle_left_transparency_texture[10][54] = 0;	doodle_left_transparency_texture[10][55] = 0;	doodle_left_transparency_texture[10][56] = 0;	doodle_left_transparency_texture[10][57] = 0;	doodle_left_transparency_texture[10][58] = 0;	doodle_left_transparency_texture[10][59] = 0;	doodle_left_transparency_texture[10][60] = 0;	doodle_left_transparency_texture[10][61] = 0;	doodle_left_transparency_texture[10][62] = 0;	doodle_left_transparency_texture[10][63] = 0;	doodle_left_transparency_texture[10][64] = 0;	doodle_left_transparency_texture[10][65] = 0;	doodle_left_transparency_texture[10][66] = 0;	doodle_left_transparency_texture[10][67] = 0;	doodle_left_transparency_texture[10][68] = 1;	doodle_left_transparency_texture[10][69] = 1;	doodle_left_transparency_texture[10][70] = 1;	doodle_left_transparency_texture[10][71] = 1;	doodle_left_transparency_texture[10][72] = 1;	doodle_left_transparency_texture[10][73] = 1;	doodle_left_transparency_texture[10][74] = 1;	doodle_left_transparency_texture[10][75] = 1;	doodle_left_transparency_texture[10][76] = 1;	doodle_left_transparency_texture[10][77] = 1;	doodle_left_transparency_texture[10][78] = 1;	doodle_left_transparency_texture[10][79] = 1;	doodle_left_transparency_texture[11][0] = 1;	doodle_left_transparency_texture[11][1] = 1;	doodle_left_transparency_texture[11][2] = 1;	doodle_left_transparency_texture[11][3] = 1;	doodle_left_transparency_texture[11][4] = 1;	doodle_left_transparency_texture[11][5] = 1;	doodle_left_transparency_texture[11][6] = 1;	doodle_left_transparency_texture[11][7] = 1;	doodle_left_transparency_texture[11][8] = 1;	doodle_left_transparency_texture[11][9] = 1;	doodle_left_transparency_texture[11][10] = 1;	doodle_left_transparency_texture[11][11] = 1;	doodle_left_transparency_texture[11][12] = 1;	doodle_left_transparency_texture[11][13] = 1;	doodle_left_transparency_texture[11][14] = 1;	doodle_left_transparency_texture[11][15] = 1;	doodle_left_transparency_texture[11][16] = 1;	doodle_left_transparency_texture[11][17] = 1;	doodle_left_transparency_texture[11][18] = 1;	doodle_left_transparency_texture[11][19] = 1;	doodle_left_transparency_texture[11][20] = 1;	doodle_left_transparency_texture[11][21] = 1;	doodle_left_transparency_texture[11][22] = 1;	doodle_left_transparency_texture[11][23] = 1;	doodle_left_transparency_texture[11][24] = 1;	doodle_left_transparency_texture[11][25] = 1;	doodle_left_transparency_texture[11][26] = 1;	doodle_left_transparency_texture[11][27] = 1;	doodle_left_transparency_texture[11][28] = 1;	doodle_left_transparency_texture[11][29] = 1;	doodle_left_transparency_texture[11][30] = 1;	doodle_left_transparency_texture[11][31] = 1;	doodle_left_transparency_texture[11][32] = 1;	doodle_left_transparency_texture[11][33] = 1;	doodle_left_transparency_texture[11][34] = 1;	doodle_left_transparency_texture[11][35] = 1;	doodle_left_transparency_texture[11][36] = 0;	doodle_left_transparency_texture[11][37] = 0;	doodle_left_transparency_texture[11][38] = 0;	doodle_left_transparency_texture[11][39] = 0;	doodle_left_transparency_texture[11][40] = 0;	doodle_left_transparency_texture[11][41] = 0;	doodle_left_transparency_texture[11][42] = 0;	doodle_left_transparency_texture[11][43] = 0;	doodle_left_transparency_texture[11][44] = 0;	doodle_left_transparency_texture[11][45] = 0;	doodle_left_transparency_texture[11][46] = 0;	doodle_left_transparency_texture[11][47] = 0;	doodle_left_transparency_texture[11][48] = 0;	doodle_left_transparency_texture[11][49] = 0;	doodle_left_transparency_texture[11][50] = 0;	doodle_left_transparency_texture[11][51] = 0;	doodle_left_transparency_texture[11][52] = 0;	doodle_left_transparency_texture[11][53] = 0;	doodle_left_transparency_texture[11][54] = 0;	doodle_left_transparency_texture[11][55] = 0;	doodle_left_transparency_texture[11][56] = 0;	doodle_left_transparency_texture[11][57] = 0;	doodle_left_transparency_texture[11][58] = 0;	doodle_left_transparency_texture[11][59] = 0;	doodle_left_transparency_texture[11][60] = 0;	doodle_left_transparency_texture[11][61] = 0;	doodle_left_transparency_texture[11][62] = 0;	doodle_left_transparency_texture[11][63] = 0;	doodle_left_transparency_texture[11][64] = 0;	doodle_left_transparency_texture[11][65] = 0;	doodle_left_transparency_texture[11][66] = 0;	doodle_left_transparency_texture[11][67] = 0;	doodle_left_transparency_texture[11][68] = 1;	doodle_left_transparency_texture[11][69] = 1;	doodle_left_transparency_texture[11][70] = 1;	doodle_left_transparency_texture[11][71] = 1;	doodle_left_transparency_texture[11][72] = 1;	doodle_left_transparency_texture[11][73] = 1;	doodle_left_transparency_texture[11][74] = 1;	doodle_left_transparency_texture[11][75] = 1;	doodle_left_transparency_texture[11][76] = 1;	doodle_left_transparency_texture[11][77] = 1;	doodle_left_transparency_texture[11][78] = 1;	doodle_left_transparency_texture[11][79] = 1;	doodle_left_transparency_texture[12][0] = 1;	doodle_left_transparency_texture[12][1] = 1;	doodle_left_transparency_texture[12][2] = 1;	doodle_left_transparency_texture[12][3] = 1;	doodle_left_transparency_texture[12][4] = 1;	doodle_left_transparency_texture[12][5] = 1;	doodle_left_transparency_texture[12][6] = 1;	doodle_left_transparency_texture[12][7] = 1;	doodle_left_transparency_texture[12][8] = 1;	doodle_left_transparency_texture[12][9] = 1;	doodle_left_transparency_texture[12][10] = 1;	doodle_left_transparency_texture[12][11] = 1;	doodle_left_transparency_texture[12][12] = 1;	doodle_left_transparency_texture[12][13] = 1;	doodle_left_transparency_texture[12][14] = 1;	doodle_left_transparency_texture[12][15] = 1;	doodle_left_transparency_texture[12][16] = 1;	doodle_left_transparency_texture[12][17] = 1;	doodle_left_transparency_texture[12][18] = 1;	doodle_left_transparency_texture[12][19] = 1;	doodle_left_transparency_texture[12][20] = 1;	doodle_left_transparency_texture[12][21] = 1;	doodle_left_transparency_texture[12][22] = 1;	doodle_left_transparency_texture[12][23] = 1;	doodle_left_transparency_texture[12][24] = 1;	doodle_left_transparency_texture[12][25] = 1;	doodle_left_transparency_texture[12][26] = 1;	doodle_left_transparency_texture[12][27] = 1;	doodle_left_transparency_texture[12][28] = 1;	doodle_left_transparency_texture[12][29] = 1;	doodle_left_transparency_texture[12][30] = 1;	doodle_left_transparency_texture[12][31] = 1;	doodle_left_transparency_texture[12][32] = 0;	doodle_left_transparency_texture[12][33] = 0;	doodle_left_transparency_texture[12][34] = 0;	doodle_left_transparency_texture[12][35] = 0;	doodle_left_transparency_texture[12][36] = 0;	doodle_left_transparency_texture[12][37] = 0;	doodle_left_transparency_texture[12][38] = 0;	doodle_left_transparency_texture[12][39] = 0;	doodle_left_transparency_texture[12][40] = 0;	doodle_left_transparency_texture[12][41] = 0;	doodle_left_transparency_texture[12][42] = 0;	doodle_left_transparency_texture[12][43] = 0;	doodle_left_transparency_texture[12][44] = 0;	doodle_left_transparency_texture[12][45] = 0;	doodle_left_transparency_texture[12][46] = 0;	doodle_left_transparency_texture[12][47] = 0;	doodle_left_transparency_texture[12][48] = 0;	doodle_left_transparency_texture[12][49] = 0;	doodle_left_transparency_texture[12][50] = 0;	doodle_left_transparency_texture[12][51] = 0;	doodle_left_transparency_texture[12][52] = 0;	doodle_left_transparency_texture[12][53] = 0;	doodle_left_transparency_texture[12][54] = 0;	doodle_left_transparency_texture[12][55] = 0;	doodle_left_transparency_texture[12][56] = 0;	doodle_left_transparency_texture[12][57] = 0;	doodle_left_transparency_texture[12][58] = 0;	doodle_left_transparency_texture[12][59] = 0;	doodle_left_transparency_texture[12][60] = 0;	doodle_left_transparency_texture[12][61] = 0;	doodle_left_transparency_texture[12][62] = 0;	doodle_left_transparency_texture[12][63] = 0;	doodle_left_transparency_texture[12][64] = 0;	doodle_left_transparency_texture[12][65] = 0;	doodle_left_transparency_texture[12][66] = 0;	doodle_left_transparency_texture[12][67] = 0;	doodle_left_transparency_texture[12][68] = 0;	doodle_left_transparency_texture[12][69] = 0;	doodle_left_transparency_texture[12][70] = 0;	doodle_left_transparency_texture[12][71] = 0;	doodle_left_transparency_texture[12][72] = 1;	doodle_left_transparency_texture[12][73] = 1;	doodle_left_transparency_texture[12][74] = 1;	doodle_left_transparency_texture[12][75] = 1;	doodle_left_transparency_texture[12][76] = 1;	doodle_left_transparency_texture[12][77] = 1;	doodle_left_transparency_texture[12][78] = 1;	doodle_left_transparency_texture[12][79] = 1;	doodle_left_transparency_texture[13][0] = 1;	doodle_left_transparency_texture[13][1] = 1;	doodle_left_transparency_texture[13][2] = 1;	doodle_left_transparency_texture[13][3] = 1;	doodle_left_transparency_texture[13][4] = 1;	doodle_left_transparency_texture[13][5] = 1;	doodle_left_transparency_texture[13][6] = 1;	doodle_left_transparency_texture[13][7] = 1;	doodle_left_transparency_texture[13][8] = 1;	doodle_left_transparency_texture[13][9] = 1;	doodle_left_transparency_texture[13][10] = 1;	doodle_left_transparency_texture[13][11] = 1;	doodle_left_transparency_texture[13][12] = 1;	doodle_left_transparency_texture[13][13] = 1;	doodle_left_transparency_texture[13][14] = 1;	doodle_left_transparency_texture[13][15] = 1;	doodle_left_transparency_texture[13][16] = 1;	doodle_left_transparency_texture[13][17] = 1;	doodle_left_transparency_texture[13][18] = 1;	doodle_left_transparency_texture[13][19] = 1;	doodle_left_transparency_texture[13][20] = 1;	doodle_left_transparency_texture[13][21] = 1;	doodle_left_transparency_texture[13][22] = 1;	doodle_left_transparency_texture[13][23] = 1;	doodle_left_transparency_texture[13][24] = 1;	doodle_left_transparency_texture[13][25] = 1;	doodle_left_transparency_texture[13][26] = 1;	doodle_left_transparency_texture[13][27] = 1;	doodle_left_transparency_texture[13][28] = 1;	doodle_left_transparency_texture[13][29] = 1;	doodle_left_transparency_texture[13][30] = 1;	doodle_left_transparency_texture[13][31] = 1;	doodle_left_transparency_texture[13][32] = 0;	doodle_left_transparency_texture[13][33] = 0;	doodle_left_transparency_texture[13][34] = 0;	doodle_left_transparency_texture[13][35] = 0;	doodle_left_transparency_texture[13][36] = 0;	doodle_left_transparency_texture[13][37] = 0;	doodle_left_transparency_texture[13][38] = 0;	doodle_left_transparency_texture[13][39] = 0;	doodle_left_transparency_texture[13][40] = 0;	doodle_left_transparency_texture[13][41] = 0;	doodle_left_transparency_texture[13][42] = 0;	doodle_left_transparency_texture[13][43] = 0;	doodle_left_transparency_texture[13][44] = 0;	doodle_left_transparency_texture[13][45] = 0;	doodle_left_transparency_texture[13][46] = 0;	doodle_left_transparency_texture[13][47] = 0;	doodle_left_transparency_texture[13][48] = 0;	doodle_left_transparency_texture[13][49] = 0;	doodle_left_transparency_texture[13][50] = 0;	doodle_left_transparency_texture[13][51] = 0;	doodle_left_transparency_texture[13][52] = 0;	doodle_left_transparency_texture[13][53] = 0;	doodle_left_transparency_texture[13][54] = 0;	doodle_left_transparency_texture[13][55] = 0;	doodle_left_transparency_texture[13][56] = 0;	doodle_left_transparency_texture[13][57] = 0;	doodle_left_transparency_texture[13][58] = 0;	doodle_left_transparency_texture[13][59] = 0;	doodle_left_transparency_texture[13][60] = 0;	doodle_left_transparency_texture[13][61] = 0;	doodle_left_transparency_texture[13][62] = 0;	doodle_left_transparency_texture[13][63] = 0;	doodle_left_transparency_texture[13][64] = 0;	doodle_left_transparency_texture[13][65] = 0;	doodle_left_transparency_texture[13][66] = 0;	doodle_left_transparency_texture[13][67] = 0;	doodle_left_transparency_texture[13][68] = 0;	doodle_left_transparency_texture[13][69] = 0;	doodle_left_transparency_texture[13][70] = 0;	doodle_left_transparency_texture[13][71] = 0;	doodle_left_transparency_texture[13][72] = 1;	doodle_left_transparency_texture[13][73] = 1;	doodle_left_transparency_texture[13][74] = 1;	doodle_left_transparency_texture[13][75] = 1;	doodle_left_transparency_texture[13][76] = 1;	doodle_left_transparency_texture[13][77] = 1;	doodle_left_transparency_texture[13][78] = 1;	doodle_left_transparency_texture[13][79] = 1;	doodle_left_transparency_texture[14][0] = 1;	doodle_left_transparency_texture[14][1] = 1;	doodle_left_transparency_texture[14][2] = 1;	doodle_left_transparency_texture[14][3] = 1;	doodle_left_transparency_texture[14][4] = 1;	doodle_left_transparency_texture[14][5] = 1;	doodle_left_transparency_texture[14][6] = 1;	doodle_left_transparency_texture[14][7] = 1;	doodle_left_transparency_texture[14][8] = 1;	doodle_left_transparency_texture[14][9] = 1;	doodle_left_transparency_texture[14][10] = 1;	doodle_left_transparency_texture[14][11] = 1;	doodle_left_transparency_texture[14][12] = 1;	doodle_left_transparency_texture[14][13] = 1;	doodle_left_transparency_texture[14][14] = 1;	doodle_left_transparency_texture[14][15] = 1;	doodle_left_transparency_texture[14][16] = 1;	doodle_left_transparency_texture[14][17] = 1;	doodle_left_transparency_texture[14][18] = 1;	doodle_left_transparency_texture[14][19] = 1;	doodle_left_transparency_texture[14][20] = 1;	doodle_left_transparency_texture[14][21] = 1;	doodle_left_transparency_texture[14][22] = 1;	doodle_left_transparency_texture[14][23] = 1;	doodle_left_transparency_texture[14][24] = 1;	doodle_left_transparency_texture[14][25] = 1;	doodle_left_transparency_texture[14][26] = 1;	doodle_left_transparency_texture[14][27] = 1;	doodle_left_transparency_texture[14][28] = 1;	doodle_left_transparency_texture[14][29] = 1;	doodle_left_transparency_texture[14][30] = 1;	doodle_left_transparency_texture[14][31] = 1;	doodle_left_transparency_texture[14][32] = 0;	doodle_left_transparency_texture[14][33] = 0;	doodle_left_transparency_texture[14][34] = 0;	doodle_left_transparency_texture[14][35] = 0;	doodle_left_transparency_texture[14][36] = 0;	doodle_left_transparency_texture[14][37] = 0;	doodle_left_transparency_texture[14][38] = 0;	doodle_left_transparency_texture[14][39] = 0;	doodle_left_transparency_texture[14][40] = 0;	doodle_left_transparency_texture[14][41] = 0;	doodle_left_transparency_texture[14][42] = 0;	doodle_left_transparency_texture[14][43] = 0;	doodle_left_transparency_texture[14][44] = 0;	doodle_left_transparency_texture[14][45] = 0;	doodle_left_transparency_texture[14][46] = 0;	doodle_left_transparency_texture[14][47] = 0;	doodle_left_transparency_texture[14][48] = 0;	doodle_left_transparency_texture[14][49] = 0;	doodle_left_transparency_texture[14][50] = 0;	doodle_left_transparency_texture[14][51] = 0;	doodle_left_transparency_texture[14][52] = 0;	doodle_left_transparency_texture[14][53] = 0;	doodle_left_transparency_texture[14][54] = 0;	doodle_left_transparency_texture[14][55] = 0;	doodle_left_transparency_texture[14][56] = 0;	doodle_left_transparency_texture[14][57] = 0;	doodle_left_transparency_texture[14][58] = 0;	doodle_left_transparency_texture[14][59] = 0;	doodle_left_transparency_texture[14][60] = 0;	doodle_left_transparency_texture[14][61] = 0;	doodle_left_transparency_texture[14][62] = 0;	doodle_left_transparency_texture[14][63] = 0;	doodle_left_transparency_texture[14][64] = 0;	doodle_left_transparency_texture[14][65] = 0;	doodle_left_transparency_texture[14][66] = 0;	doodle_left_transparency_texture[14][67] = 0;	doodle_left_transparency_texture[14][68] = 0;	doodle_left_transparency_texture[14][69] = 0;	doodle_left_transparency_texture[14][70] = 0;	doodle_left_transparency_texture[14][71] = 0;	doodle_left_transparency_texture[14][72] = 1;	doodle_left_transparency_texture[14][73] = 1;	doodle_left_transparency_texture[14][74] = 1;	doodle_left_transparency_texture[14][75] = 1;	doodle_left_transparency_texture[14][76] = 1;	doodle_left_transparency_texture[14][77] = 1;	doodle_left_transparency_texture[14][78] = 1;	doodle_left_transparency_texture[14][79] = 1;	doodle_left_transparency_texture[15][0] = 1;	doodle_left_transparency_texture[15][1] = 1;	doodle_left_transparency_texture[15][2] = 1;	doodle_left_transparency_texture[15][3] = 1;	doodle_left_transparency_texture[15][4] = 1;	doodle_left_transparency_texture[15][5] = 1;	doodle_left_transparency_texture[15][6] = 1;	doodle_left_transparency_texture[15][7] = 1;	doodle_left_transparency_texture[15][8] = 1;	doodle_left_transparency_texture[15][9] = 1;	doodle_left_transparency_texture[15][10] = 1;	doodle_left_transparency_texture[15][11] = 1;	doodle_left_transparency_texture[15][12] = 1;	doodle_left_transparency_texture[15][13] = 1;	doodle_left_transparency_texture[15][14] = 1;	doodle_left_transparency_texture[15][15] = 1;	doodle_left_transparency_texture[15][16] = 1;	doodle_left_transparency_texture[15][17] = 1;	doodle_left_transparency_texture[15][18] = 1;	doodle_left_transparency_texture[15][19] = 1;	doodle_left_transparency_texture[15][20] = 1;	doodle_left_transparency_texture[15][21] = 1;	doodle_left_transparency_texture[15][22] = 1;	doodle_left_transparency_texture[15][23] = 1;	doodle_left_transparency_texture[15][24] = 1;	doodle_left_transparency_texture[15][25] = 1;	doodle_left_transparency_texture[15][26] = 1;	doodle_left_transparency_texture[15][27] = 1;	doodle_left_transparency_texture[15][28] = 1;	doodle_left_transparency_texture[15][29] = 1;	doodle_left_transparency_texture[15][30] = 1;	doodle_left_transparency_texture[15][31] = 1;	doodle_left_transparency_texture[15][32] = 0;	doodle_left_transparency_texture[15][33] = 0;	doodle_left_transparency_texture[15][34] = 0;	doodle_left_transparency_texture[15][35] = 0;	doodle_left_transparency_texture[15][36] = 0;	doodle_left_transparency_texture[15][37] = 0;	doodle_left_transparency_texture[15][38] = 0;	doodle_left_transparency_texture[15][39] = 0;	doodle_left_transparency_texture[15][40] = 0;	doodle_left_transparency_texture[15][41] = 0;	doodle_left_transparency_texture[15][42] = 0;	doodle_left_transparency_texture[15][43] = 0;	doodle_left_transparency_texture[15][44] = 0;	doodle_left_transparency_texture[15][45] = 0;	doodle_left_transparency_texture[15][46] = 0;	doodle_left_transparency_texture[15][47] = 0;	doodle_left_transparency_texture[15][48] = 0;	doodle_left_transparency_texture[15][49] = 0;	doodle_left_transparency_texture[15][50] = 0;	doodle_left_transparency_texture[15][51] = 0;	doodle_left_transparency_texture[15][52] = 0;	doodle_left_transparency_texture[15][53] = 0;	doodle_left_transparency_texture[15][54] = 0;	doodle_left_transparency_texture[15][55] = 0;	doodle_left_transparency_texture[15][56] = 0;	doodle_left_transparency_texture[15][57] = 0;	doodle_left_transparency_texture[15][58] = 0;	doodle_left_transparency_texture[15][59] = 0;	doodle_left_transparency_texture[15][60] = 0;	doodle_left_transparency_texture[15][61] = 0;	doodle_left_transparency_texture[15][62] = 0;	doodle_left_transparency_texture[15][63] = 0;	doodle_left_transparency_texture[15][64] = 0;	doodle_left_transparency_texture[15][65] = 0;	doodle_left_transparency_texture[15][66] = 0;	doodle_left_transparency_texture[15][67] = 0;	doodle_left_transparency_texture[15][68] = 0;	doodle_left_transparency_texture[15][69] = 0;	doodle_left_transparency_texture[15][70] = 0;	doodle_left_transparency_texture[15][71] = 0;	doodle_left_transparency_texture[15][72] = 1;	doodle_left_transparency_texture[15][73] = 1;	doodle_left_transparency_texture[15][74] = 1;	doodle_left_transparency_texture[15][75] = 1;	doodle_left_transparency_texture[15][76] = 1;	doodle_left_transparency_texture[15][77] = 1;	doodle_left_transparency_texture[15][78] = 1;	doodle_left_transparency_texture[15][79] = 1;	doodle_left_transparency_texture[16][0] = 1;	doodle_left_transparency_texture[16][1] = 1;	doodle_left_transparency_texture[16][2] = 1;	doodle_left_transparency_texture[16][3] = 1;	doodle_left_transparency_texture[16][4] = 1;	doodle_left_transparency_texture[16][5] = 1;	doodle_left_transparency_texture[16][6] = 1;	doodle_left_transparency_texture[16][7] = 1;	doodle_left_transparency_texture[16][8] = 1;	doodle_left_transparency_texture[16][9] = 1;	doodle_left_transparency_texture[16][10] = 1;	doodle_left_transparency_texture[16][11] = 1;	doodle_left_transparency_texture[16][12] = 1;	doodle_left_transparency_texture[16][13] = 1;	doodle_left_transparency_texture[16][14] = 1;	doodle_left_transparency_texture[16][15] = 1;	doodle_left_transparency_texture[16][16] = 1;	doodle_left_transparency_texture[16][17] = 1;	doodle_left_transparency_texture[16][18] = 1;	doodle_left_transparency_texture[16][19] = 1;	doodle_left_transparency_texture[16][20] = 1;	doodle_left_transparency_texture[16][21] = 1;	doodle_left_transparency_texture[16][22] = 1;	doodle_left_transparency_texture[16][23] = 1;	doodle_left_transparency_texture[16][24] = 1;	doodle_left_transparency_texture[16][25] = 1;	doodle_left_transparency_texture[16][26] = 1;	doodle_left_transparency_texture[16][27] = 1;	doodle_left_transparency_texture[16][28] = 0;	doodle_left_transparency_texture[16][29] = 0;	doodle_left_transparency_texture[16][30] = 0;	doodle_left_transparency_texture[16][31] = 0;	doodle_left_transparency_texture[16][32] = 0;	doodle_left_transparency_texture[16][33] = 0;	doodle_left_transparency_texture[16][34] = 0;	doodle_left_transparency_texture[16][35] = 0;	doodle_left_transparency_texture[16][36] = 0;	doodle_left_transparency_texture[16][37] = 0;	doodle_left_transparency_texture[16][38] = 0;	doodle_left_transparency_texture[16][39] = 0;	doodle_left_transparency_texture[16][40] = 0;	doodle_left_transparency_texture[16][41] = 0;	doodle_left_transparency_texture[16][42] = 0;	doodle_left_transparency_texture[16][43] = 0;	doodle_left_transparency_texture[16][44] = 0;	doodle_left_transparency_texture[16][45] = 0;	doodle_left_transparency_texture[16][46] = 0;	doodle_left_transparency_texture[16][47] = 0;	doodle_left_transparency_texture[16][48] = 0;	doodle_left_transparency_texture[16][49] = 0;	doodle_left_transparency_texture[16][50] = 0;	doodle_left_transparency_texture[16][51] = 0;	doodle_left_transparency_texture[16][52] = 0;	doodle_left_transparency_texture[16][53] = 0;	doodle_left_transparency_texture[16][54] = 0;	doodle_left_transparency_texture[16][55] = 0;	doodle_left_transparency_texture[16][56] = 0;	doodle_left_transparency_texture[16][57] = 0;	doodle_left_transparency_texture[16][58] = 0;	doodle_left_transparency_texture[16][59] = 0;	doodle_left_transparency_texture[16][60] = 0;	doodle_left_transparency_texture[16][61] = 0;	doodle_left_transparency_texture[16][62] = 0;	doodle_left_transparency_texture[16][63] = 0;	doodle_left_transparency_texture[16][64] = 0;	doodle_left_transparency_texture[16][65] = 0;	doodle_left_transparency_texture[16][66] = 0;	doodle_left_transparency_texture[16][67] = 0;	doodle_left_transparency_texture[16][68] = 0;	doodle_left_transparency_texture[16][69] = 0;	doodle_left_transparency_texture[16][70] = 0;	doodle_left_transparency_texture[16][71] = 0;	doodle_left_transparency_texture[16][72] = 0;	doodle_left_transparency_texture[16][73] = 0;	doodle_left_transparency_texture[16][74] = 0;	doodle_left_transparency_texture[16][75] = 0;	doodle_left_transparency_texture[16][76] = 1;	doodle_left_transparency_texture[16][77] = 1;	doodle_left_transparency_texture[16][78] = 1;	doodle_left_transparency_texture[16][79] = 1;	doodle_left_transparency_texture[17][0] = 1;	doodle_left_transparency_texture[17][1] = 1;	doodle_left_transparency_texture[17][2] = 1;	doodle_left_transparency_texture[17][3] = 1;	doodle_left_transparency_texture[17][4] = 1;	doodle_left_transparency_texture[17][5] = 1;	doodle_left_transparency_texture[17][6] = 1;	doodle_left_transparency_texture[17][7] = 1;	doodle_left_transparency_texture[17][8] = 1;	doodle_left_transparency_texture[17][9] = 1;	doodle_left_transparency_texture[17][10] = 1;	doodle_left_transparency_texture[17][11] = 1;	doodle_left_transparency_texture[17][12] = 1;	doodle_left_transparency_texture[17][13] = 1;	doodle_left_transparency_texture[17][14] = 1;	doodle_left_transparency_texture[17][15] = 1;	doodle_left_transparency_texture[17][16] = 1;	doodle_left_transparency_texture[17][17] = 1;	doodle_left_transparency_texture[17][18] = 1;	doodle_left_transparency_texture[17][19] = 1;	doodle_left_transparency_texture[17][20] = 1;	doodle_left_transparency_texture[17][21] = 1;	doodle_left_transparency_texture[17][22] = 1;	doodle_left_transparency_texture[17][23] = 1;	doodle_left_transparency_texture[17][24] = 1;	doodle_left_transparency_texture[17][25] = 1;	doodle_left_transparency_texture[17][26] = 1;	doodle_left_transparency_texture[17][27] = 1;	doodle_left_transparency_texture[17][28] = 0;	doodle_left_transparency_texture[17][29] = 0;	doodle_left_transparency_texture[17][30] = 0;	doodle_left_transparency_texture[17][31] = 0;	doodle_left_transparency_texture[17][32] = 0;	doodle_left_transparency_texture[17][33] = 0;	doodle_left_transparency_texture[17][34] = 0;	doodle_left_transparency_texture[17][35] = 0;	doodle_left_transparency_texture[17][36] = 0;	doodle_left_transparency_texture[17][37] = 0;	doodle_left_transparency_texture[17][38] = 0;	doodle_left_transparency_texture[17][39] = 0;	doodle_left_transparency_texture[17][40] = 0;	doodle_left_transparency_texture[17][41] = 0;	doodle_left_transparency_texture[17][42] = 0;	doodle_left_transparency_texture[17][43] = 0;	doodle_left_transparency_texture[17][44] = 0;	doodle_left_transparency_texture[17][45] = 0;	doodle_left_transparency_texture[17][46] = 0;	doodle_left_transparency_texture[17][47] = 0;	doodle_left_transparency_texture[17][48] = 0;	doodle_left_transparency_texture[17][49] = 0;	doodle_left_transparency_texture[17][50] = 0;	doodle_left_transparency_texture[17][51] = 0;	doodle_left_transparency_texture[17][52] = 0;	doodle_left_transparency_texture[17][53] = 0;	doodle_left_transparency_texture[17][54] = 0;	doodle_left_transparency_texture[17][55] = 0;	doodle_left_transparency_texture[17][56] = 0;	doodle_left_transparency_texture[17][57] = 0;	doodle_left_transparency_texture[17][58] = 0;	doodle_left_transparency_texture[17][59] = 0;	doodle_left_transparency_texture[17][60] = 0;	doodle_left_transparency_texture[17][61] = 0;	doodle_left_transparency_texture[17][62] = 0;	doodle_left_transparency_texture[17][63] = 0;	doodle_left_transparency_texture[17][64] = 0;	doodle_left_transparency_texture[17][65] = 0;	doodle_left_transparency_texture[17][66] = 0;	doodle_left_transparency_texture[17][67] = 0;	doodle_left_transparency_texture[17][68] = 0;	doodle_left_transparency_texture[17][69] = 0;	doodle_left_transparency_texture[17][70] = 0;	doodle_left_transparency_texture[17][71] = 0;	doodle_left_transparency_texture[17][72] = 0;	doodle_left_transparency_texture[17][73] = 0;	doodle_left_transparency_texture[17][74] = 0;	doodle_left_transparency_texture[17][75] = 0;	doodle_left_transparency_texture[17][76] = 1;	doodle_left_transparency_texture[17][77] = 1;	doodle_left_transparency_texture[17][78] = 1;	doodle_left_transparency_texture[17][79] = 1;	doodle_left_transparency_texture[18][0] = 1;	doodle_left_transparency_texture[18][1] = 1;	doodle_left_transparency_texture[18][2] = 1;	doodle_left_transparency_texture[18][3] = 1;	doodle_left_transparency_texture[18][4] = 1;	doodle_left_transparency_texture[18][5] = 1;	doodle_left_transparency_texture[18][6] = 1;	doodle_left_transparency_texture[18][7] = 1;	doodle_left_transparency_texture[18][8] = 1;	doodle_left_transparency_texture[18][9] = 1;	doodle_left_transparency_texture[18][10] = 1;	doodle_left_transparency_texture[18][11] = 1;	doodle_left_transparency_texture[18][12] = 1;	doodle_left_transparency_texture[18][13] = 1;	doodle_left_transparency_texture[18][14] = 1;	doodle_left_transparency_texture[18][15] = 1;	doodle_left_transparency_texture[18][16] = 1;	doodle_left_transparency_texture[18][17] = 1;	doodle_left_transparency_texture[18][18] = 1;	doodle_left_transparency_texture[18][19] = 1;	doodle_left_transparency_texture[18][20] = 1;	doodle_left_transparency_texture[18][21] = 1;	doodle_left_transparency_texture[18][22] = 1;	doodle_left_transparency_texture[18][23] = 1;	doodle_left_transparency_texture[18][24] = 1;	doodle_left_transparency_texture[18][25] = 1;	doodle_left_transparency_texture[18][26] = 1;	doodle_left_transparency_texture[18][27] = 1;	doodle_left_transparency_texture[18][28] = 0;	doodle_left_transparency_texture[18][29] = 0;	doodle_left_transparency_texture[18][30] = 0;	doodle_left_transparency_texture[18][31] = 0;	doodle_left_transparency_texture[18][32] = 0;	doodle_left_transparency_texture[18][33] = 0;	doodle_left_transparency_texture[18][34] = 0;	doodle_left_transparency_texture[18][35] = 0;	doodle_left_transparency_texture[18][36] = 0;	doodle_left_transparency_texture[18][37] = 0;	doodle_left_transparency_texture[18][38] = 0;	doodle_left_transparency_texture[18][39] = 0;	doodle_left_transparency_texture[18][40] = 0;	doodle_left_transparency_texture[18][41] = 0;	doodle_left_transparency_texture[18][42] = 0;	doodle_left_transparency_texture[18][43] = 0;	doodle_left_transparency_texture[18][44] = 0;	doodle_left_transparency_texture[18][45] = 0;	doodle_left_transparency_texture[18][46] = 0;	doodle_left_transparency_texture[18][47] = 0;	doodle_left_transparency_texture[18][48] = 0;	doodle_left_transparency_texture[18][49] = 0;	doodle_left_transparency_texture[18][50] = 0;	doodle_left_transparency_texture[18][51] = 0;	doodle_left_transparency_texture[18][52] = 0;	doodle_left_transparency_texture[18][53] = 0;	doodle_left_transparency_texture[18][54] = 0;	doodle_left_transparency_texture[18][55] = 0;	doodle_left_transparency_texture[18][56] = 0;	doodle_left_transparency_texture[18][57] = 0;	doodle_left_transparency_texture[18][58] = 0;	doodle_left_transparency_texture[18][59] = 0;	doodle_left_transparency_texture[18][60] = 0;	doodle_left_transparency_texture[18][61] = 0;	doodle_left_transparency_texture[18][62] = 0;	doodle_left_transparency_texture[18][63] = 0;	doodle_left_transparency_texture[18][64] = 0;	doodle_left_transparency_texture[18][65] = 0;	doodle_left_transparency_texture[18][66] = 0;	doodle_left_transparency_texture[18][67] = 0;	doodle_left_transparency_texture[18][68] = 0;	doodle_left_transparency_texture[18][69] = 0;	doodle_left_transparency_texture[18][70] = 0;	doodle_left_transparency_texture[18][71] = 0;	doodle_left_transparency_texture[18][72] = 0;	doodle_left_transparency_texture[18][73] = 0;	doodle_left_transparency_texture[18][74] = 0;	doodle_left_transparency_texture[18][75] = 0;	doodle_left_transparency_texture[18][76] = 1;	doodle_left_transparency_texture[18][77] = 1;	doodle_left_transparency_texture[18][78] = 1;	doodle_left_transparency_texture[18][79] = 1;	doodle_left_transparency_texture[19][0] = 1;	doodle_left_transparency_texture[19][1] = 1;	doodle_left_transparency_texture[19][2] = 1;	doodle_left_transparency_texture[19][3] = 1;	doodle_left_transparency_texture[19][4] = 1;	doodle_left_transparency_texture[19][5] = 1;	doodle_left_transparency_texture[19][6] = 1;	doodle_left_transparency_texture[19][7] = 1;	doodle_left_transparency_texture[19][8] = 1;	doodle_left_transparency_texture[19][9] = 1;	doodle_left_transparency_texture[19][10] = 1;	doodle_left_transparency_texture[19][11] = 1;	doodle_left_transparency_texture[19][12] = 1;	doodle_left_transparency_texture[19][13] = 1;	doodle_left_transparency_texture[19][14] = 1;	doodle_left_transparency_texture[19][15] = 1;	doodle_left_transparency_texture[19][16] = 1;	doodle_left_transparency_texture[19][17] = 1;	doodle_left_transparency_texture[19][18] = 1;	doodle_left_transparency_texture[19][19] = 1;	doodle_left_transparency_texture[19][20] = 1;	doodle_left_transparency_texture[19][21] = 1;	doodle_left_transparency_texture[19][22] = 1;	doodle_left_transparency_texture[19][23] = 1;	doodle_left_transparency_texture[19][24] = 1;	doodle_left_transparency_texture[19][25] = 1;	doodle_left_transparency_texture[19][26] = 1;	doodle_left_transparency_texture[19][27] = 1;	doodle_left_transparency_texture[19][28] = 0;	doodle_left_transparency_texture[19][29] = 0;	doodle_left_transparency_texture[19][30] = 0;	doodle_left_transparency_texture[19][31] = 0;	doodle_left_transparency_texture[19][32] = 0;	doodle_left_transparency_texture[19][33] = 0;	doodle_left_transparency_texture[19][34] = 0;	doodle_left_transparency_texture[19][35] = 0;	doodle_left_transparency_texture[19][36] = 0;	doodle_left_transparency_texture[19][37] = 0;	doodle_left_transparency_texture[19][38] = 0;	doodle_left_transparency_texture[19][39] = 0;	doodle_left_transparency_texture[19][40] = 0;	doodle_left_transparency_texture[19][41] = 0;	doodle_left_transparency_texture[19][42] = 0;	doodle_left_transparency_texture[19][43] = 0;	doodle_left_transparency_texture[19][44] = 0;	doodle_left_transparency_texture[19][45] = 0;	doodle_left_transparency_texture[19][46] = 0;	doodle_left_transparency_texture[19][47] = 0;	doodle_left_transparency_texture[19][48] = 0;	doodle_left_transparency_texture[19][49] = 0;	doodle_left_transparency_texture[19][50] = 0;	doodle_left_transparency_texture[19][51] = 0;	doodle_left_transparency_texture[19][52] = 0;	doodle_left_transparency_texture[19][53] = 0;	doodle_left_transparency_texture[19][54] = 0;	doodle_left_transparency_texture[19][55] = 0;	doodle_left_transparency_texture[19][56] = 0;	doodle_left_transparency_texture[19][57] = 0;	doodle_left_transparency_texture[19][58] = 0;	doodle_left_transparency_texture[19][59] = 0;	doodle_left_transparency_texture[19][60] = 0;	doodle_left_transparency_texture[19][61] = 0;	doodle_left_transparency_texture[19][62] = 0;	doodle_left_transparency_texture[19][63] = 0;	doodle_left_transparency_texture[19][64] = 0;	doodle_left_transparency_texture[19][65] = 0;	doodle_left_transparency_texture[19][66] = 0;	doodle_left_transparency_texture[19][67] = 0;	doodle_left_transparency_texture[19][68] = 0;	doodle_left_transparency_texture[19][69] = 0;	doodle_left_transparency_texture[19][70] = 0;	doodle_left_transparency_texture[19][71] = 0;	doodle_left_transparency_texture[19][72] = 0;	doodle_left_transparency_texture[19][73] = 0;	doodle_left_transparency_texture[19][74] = 0;	doodle_left_transparency_texture[19][75] = 0;	doodle_left_transparency_texture[19][76] = 1;	doodle_left_transparency_texture[19][77] = 1;	doodle_left_transparency_texture[19][78] = 1;	doodle_left_transparency_texture[19][79] = 1;	doodle_left_transparency_texture[20][0] = 1;	doodle_left_transparency_texture[20][1] = 1;	doodle_left_transparency_texture[20][2] = 1;	doodle_left_transparency_texture[20][3] = 1;	doodle_left_transparency_texture[20][4] = 1;	doodle_left_transparency_texture[20][5] = 1;	doodle_left_transparency_texture[20][6] = 1;	doodle_left_transparency_texture[20][7] = 1;	doodle_left_transparency_texture[20][8] = 1;	doodle_left_transparency_texture[20][9] = 1;	doodle_left_transparency_texture[20][10] = 1;	doodle_left_transparency_texture[20][11] = 1;	doodle_left_transparency_texture[20][12] = 1;	doodle_left_transparency_texture[20][13] = 1;	doodle_left_transparency_texture[20][14] = 1;	doodle_left_transparency_texture[20][15] = 1;	doodle_left_transparency_texture[20][16] = 1;	doodle_left_transparency_texture[20][17] = 1;	doodle_left_transparency_texture[20][18] = 1;	doodle_left_transparency_texture[20][19] = 1;	doodle_left_transparency_texture[20][20] = 1;	doodle_left_transparency_texture[20][21] = 1;	doodle_left_transparency_texture[20][22] = 1;	doodle_left_transparency_texture[20][23] = 1;	doodle_left_transparency_texture[20][24] = 1;	doodle_left_transparency_texture[20][25] = 1;	doodle_left_transparency_texture[20][26] = 1;	doodle_left_transparency_texture[20][27] = 1;	doodle_left_transparency_texture[20][28] = 0;	doodle_left_transparency_texture[20][29] = 0;	doodle_left_transparency_texture[20][30] = 0;	doodle_left_transparency_texture[20][31] = 0;	doodle_left_transparency_texture[20][32] = 0;	doodle_left_transparency_texture[20][33] = 0;	doodle_left_transparency_texture[20][34] = 0;	doodle_left_transparency_texture[20][35] = 0;	doodle_left_transparency_texture[20][36] = 0;	doodle_left_transparency_texture[20][37] = 0;	doodle_left_transparency_texture[20][38] = 0;	doodle_left_transparency_texture[20][39] = 0;	doodle_left_transparency_texture[20][40] = 0;	doodle_left_transparency_texture[20][41] = 0;	doodle_left_transparency_texture[20][42] = 0;	doodle_left_transparency_texture[20][43] = 0;	doodle_left_transparency_texture[20][44] = 0;	doodle_left_transparency_texture[20][45] = 0;	doodle_left_transparency_texture[20][46] = 0;	doodle_left_transparency_texture[20][47] = 0;	doodle_left_transparency_texture[20][48] = 0;	doodle_left_transparency_texture[20][49] = 0;	doodle_left_transparency_texture[20][50] = 0;	doodle_left_transparency_texture[20][51] = 0;	doodle_left_transparency_texture[20][52] = 0;	doodle_left_transparency_texture[20][53] = 0;	doodle_left_transparency_texture[20][54] = 0;	doodle_left_transparency_texture[20][55] = 0;	doodle_left_transparency_texture[20][56] = 0;	doodle_left_transparency_texture[20][57] = 0;	doodle_left_transparency_texture[20][58] = 0;	doodle_left_transparency_texture[20][59] = 0;	doodle_left_transparency_texture[20][60] = 0;	doodle_left_transparency_texture[20][61] = 0;	doodle_left_transparency_texture[20][62] = 0;	doodle_left_transparency_texture[20][63] = 0;	doodle_left_transparency_texture[20][64] = 0;	doodle_left_transparency_texture[20][65] = 0;	doodle_left_transparency_texture[20][66] = 0;	doodle_left_transparency_texture[20][67] = 0;	doodle_left_transparency_texture[20][68] = 0;	doodle_left_transparency_texture[20][69] = 0;	doodle_left_transparency_texture[20][70] = 0;	doodle_left_transparency_texture[20][71] = 0;	doodle_left_transparency_texture[20][72] = 0;	doodle_left_transparency_texture[20][73] = 0;	doodle_left_transparency_texture[20][74] = 0;	doodle_left_transparency_texture[20][75] = 0;	doodle_left_transparency_texture[20][76] = 1;	doodle_left_transparency_texture[20][77] = 1;	doodle_left_transparency_texture[20][78] = 1;	doodle_left_transparency_texture[20][79] = 1;	doodle_left_transparency_texture[21][0] = 1;	doodle_left_transparency_texture[21][1] = 1;	doodle_left_transparency_texture[21][2] = 1;	doodle_left_transparency_texture[21][3] = 1;	doodle_left_transparency_texture[21][4] = 1;	doodle_left_transparency_texture[21][5] = 1;	doodle_left_transparency_texture[21][6] = 1;	doodle_left_transparency_texture[21][7] = 1;	doodle_left_transparency_texture[21][8] = 1;	doodle_left_transparency_texture[21][9] = 1;	doodle_left_transparency_texture[21][10] = 1;	doodle_left_transparency_texture[21][11] = 1;	doodle_left_transparency_texture[21][12] = 1;	doodle_left_transparency_texture[21][13] = 1;	doodle_left_transparency_texture[21][14] = 1;	doodle_left_transparency_texture[21][15] = 1;	doodle_left_transparency_texture[21][16] = 1;	doodle_left_transparency_texture[21][17] = 1;	doodle_left_transparency_texture[21][18] = 1;	doodle_left_transparency_texture[21][19] = 1;	doodle_left_transparency_texture[21][20] = 1;	doodle_left_transparency_texture[21][21] = 1;	doodle_left_transparency_texture[21][22] = 1;	doodle_left_transparency_texture[21][23] = 1;	doodle_left_transparency_texture[21][24] = 1;	doodle_left_transparency_texture[21][25] = 1;	doodle_left_transparency_texture[21][26] = 1;	doodle_left_transparency_texture[21][27] = 1;	doodle_left_transparency_texture[21][28] = 0;	doodle_left_transparency_texture[21][29] = 0;	doodle_left_transparency_texture[21][30] = 0;	doodle_left_transparency_texture[21][31] = 0;	doodle_left_transparency_texture[21][32] = 0;	doodle_left_transparency_texture[21][33] = 0;	doodle_left_transparency_texture[21][34] = 0;	doodle_left_transparency_texture[21][35] = 0;	doodle_left_transparency_texture[21][36] = 0;	doodle_left_transparency_texture[21][37] = 0;	doodle_left_transparency_texture[21][38] = 0;	doodle_left_transparency_texture[21][39] = 0;	doodle_left_transparency_texture[21][40] = 0;	doodle_left_transparency_texture[21][41] = 0;	doodle_left_transparency_texture[21][42] = 0;	doodle_left_transparency_texture[21][43] = 0;	doodle_left_transparency_texture[21][44] = 0;	doodle_left_transparency_texture[21][45] = 0;	doodle_left_transparency_texture[21][46] = 0;	doodle_left_transparency_texture[21][47] = 0;	doodle_left_transparency_texture[21][48] = 0;	doodle_left_transparency_texture[21][49] = 0;	doodle_left_transparency_texture[21][50] = 0;	doodle_left_transparency_texture[21][51] = 0;	doodle_left_transparency_texture[21][52] = 0;	doodle_left_transparency_texture[21][53] = 0;	doodle_left_transparency_texture[21][54] = 0;	doodle_left_transparency_texture[21][55] = 0;	doodle_left_transparency_texture[21][56] = 0;	doodle_left_transparency_texture[21][57] = 0;	doodle_left_transparency_texture[21][58] = 0;	doodle_left_transparency_texture[21][59] = 0;	doodle_left_transparency_texture[21][60] = 0;	doodle_left_transparency_texture[21][61] = 0;	doodle_left_transparency_texture[21][62] = 0;	doodle_left_transparency_texture[21][63] = 0;	doodle_left_transparency_texture[21][64] = 0;	doodle_left_transparency_texture[21][65] = 0;	doodle_left_transparency_texture[21][66] = 0;	doodle_left_transparency_texture[21][67] = 0;	doodle_left_transparency_texture[21][68] = 0;	doodle_left_transparency_texture[21][69] = 0;	doodle_left_transparency_texture[21][70] = 0;	doodle_left_transparency_texture[21][71] = 0;	doodle_left_transparency_texture[21][72] = 0;	doodle_left_transparency_texture[21][73] = 0;	doodle_left_transparency_texture[21][74] = 0;	doodle_left_transparency_texture[21][75] = 0;	doodle_left_transparency_texture[21][76] = 1;	doodle_left_transparency_texture[21][77] = 1;	doodle_left_transparency_texture[21][78] = 1;	doodle_left_transparency_texture[21][79] = 1;	doodle_left_transparency_texture[22][0] = 1;	doodle_left_transparency_texture[22][1] = 1;	doodle_left_transparency_texture[22][2] = 1;	doodle_left_transparency_texture[22][3] = 1;	doodle_left_transparency_texture[22][4] = 1;	doodle_left_transparency_texture[22][5] = 1;	doodle_left_transparency_texture[22][6] = 1;	doodle_left_transparency_texture[22][7] = 1;	doodle_left_transparency_texture[22][8] = 1;	doodle_left_transparency_texture[22][9] = 1;	doodle_left_transparency_texture[22][10] = 1;	doodle_left_transparency_texture[22][11] = 1;	doodle_left_transparency_texture[22][12] = 1;	doodle_left_transparency_texture[22][13] = 1;	doodle_left_transparency_texture[22][14] = 1;	doodle_left_transparency_texture[22][15] = 1;	doodle_left_transparency_texture[22][16] = 1;	doodle_left_transparency_texture[22][17] = 1;	doodle_left_transparency_texture[22][18] = 1;	doodle_left_transparency_texture[22][19] = 1;	doodle_left_transparency_texture[22][20] = 1;	doodle_left_transparency_texture[22][21] = 1;	doodle_left_transparency_texture[22][22] = 1;	doodle_left_transparency_texture[22][23] = 1;	doodle_left_transparency_texture[22][24] = 1;	doodle_left_transparency_texture[22][25] = 1;	doodle_left_transparency_texture[22][26] = 1;	doodle_left_transparency_texture[22][27] = 1;	doodle_left_transparency_texture[22][28] = 0;	doodle_left_transparency_texture[22][29] = 0;	doodle_left_transparency_texture[22][30] = 0;	doodle_left_transparency_texture[22][31] = 0;	doodle_left_transparency_texture[22][32] = 0;	doodle_left_transparency_texture[22][33] = 0;	doodle_left_transparency_texture[22][34] = 0;	doodle_left_transparency_texture[22][35] = 0;	doodle_left_transparency_texture[22][36] = 0;	doodle_left_transparency_texture[22][37] = 0;	doodle_left_transparency_texture[22][38] = 0;	doodle_left_transparency_texture[22][39] = 0;	doodle_left_transparency_texture[22][40] = 0;	doodle_left_transparency_texture[22][41] = 0;	doodle_left_transparency_texture[22][42] = 0;	doodle_left_transparency_texture[22][43] = 0;	doodle_left_transparency_texture[22][44] = 0;	doodle_left_transparency_texture[22][45] = 0;	doodle_left_transparency_texture[22][46] = 0;	doodle_left_transparency_texture[22][47] = 0;	doodle_left_transparency_texture[22][48] = 0;	doodle_left_transparency_texture[22][49] = 0;	doodle_left_transparency_texture[22][50] = 0;	doodle_left_transparency_texture[22][51] = 0;	doodle_left_transparency_texture[22][52] = 0;	doodle_left_transparency_texture[22][53] = 0;	doodle_left_transparency_texture[22][54] = 0;	doodle_left_transparency_texture[22][55] = 0;	doodle_left_transparency_texture[22][56] = 0;	doodle_left_transparency_texture[22][57] = 0;	doodle_left_transparency_texture[22][58] = 0;	doodle_left_transparency_texture[22][59] = 0;	doodle_left_transparency_texture[22][60] = 0;	doodle_left_transparency_texture[22][61] = 0;	doodle_left_transparency_texture[22][62] = 0;	doodle_left_transparency_texture[22][63] = 0;	doodle_left_transparency_texture[22][64] = 0;	doodle_left_transparency_texture[22][65] = 0;	doodle_left_transparency_texture[22][66] = 0;	doodle_left_transparency_texture[22][67] = 0;	doodle_left_transparency_texture[22][68] = 0;	doodle_left_transparency_texture[22][69] = 0;	doodle_left_transparency_texture[22][70] = 0;	doodle_left_transparency_texture[22][71] = 0;	doodle_left_transparency_texture[22][72] = 0;	doodle_left_transparency_texture[22][73] = 0;	doodle_left_transparency_texture[22][74] = 0;	doodle_left_transparency_texture[22][75] = 0;	doodle_left_transparency_texture[22][76] = 1;	doodle_left_transparency_texture[22][77] = 1;	doodle_left_transparency_texture[22][78] = 1;	doodle_left_transparency_texture[22][79] = 1;	doodle_left_transparency_texture[23][0] = 1;	doodle_left_transparency_texture[23][1] = 1;	doodle_left_transparency_texture[23][2] = 1;	doodle_left_transparency_texture[23][3] = 1;	doodle_left_transparency_texture[23][4] = 1;	doodle_left_transparency_texture[23][5] = 1;	doodle_left_transparency_texture[23][6] = 1;	doodle_left_transparency_texture[23][7] = 1;	doodle_left_transparency_texture[23][8] = 1;	doodle_left_transparency_texture[23][9] = 1;	doodle_left_transparency_texture[23][10] = 1;	doodle_left_transparency_texture[23][11] = 1;	doodle_left_transparency_texture[23][12] = 1;	doodle_left_transparency_texture[23][13] = 1;	doodle_left_transparency_texture[23][14] = 1;	doodle_left_transparency_texture[23][15] = 1;	doodle_left_transparency_texture[23][16] = 1;	doodle_left_transparency_texture[23][17] = 1;	doodle_left_transparency_texture[23][18] = 1;	doodle_left_transparency_texture[23][19] = 1;	doodle_left_transparency_texture[23][20] = 1;	doodle_left_transparency_texture[23][21] = 1;	doodle_left_transparency_texture[23][22] = 1;	doodle_left_transparency_texture[23][23] = 1;	doodle_left_transparency_texture[23][24] = 1;	doodle_left_transparency_texture[23][25] = 1;	doodle_left_transparency_texture[23][26] = 1;	doodle_left_transparency_texture[23][27] = 1;	doodle_left_transparency_texture[23][28] = 0;	doodle_left_transparency_texture[23][29] = 0;	doodle_left_transparency_texture[23][30] = 0;	doodle_left_transparency_texture[23][31] = 0;	doodle_left_transparency_texture[23][32] = 0;	doodle_left_transparency_texture[23][33] = 0;	doodle_left_transparency_texture[23][34] = 0;	doodle_left_transparency_texture[23][35] = 0;	doodle_left_transparency_texture[23][36] = 0;	doodle_left_transparency_texture[23][37] = 0;	doodle_left_transparency_texture[23][38] = 0;	doodle_left_transparency_texture[23][39] = 0;	doodle_left_transparency_texture[23][40] = 0;	doodle_left_transparency_texture[23][41] = 0;	doodle_left_transparency_texture[23][42] = 0;	doodle_left_transparency_texture[23][43] = 0;	doodle_left_transparency_texture[23][44] = 0;	doodle_left_transparency_texture[23][45] = 0;	doodle_left_transparency_texture[23][46] = 0;	doodle_left_transparency_texture[23][47] = 0;	doodle_left_transparency_texture[23][48] = 0;	doodle_left_transparency_texture[23][49] = 0;	doodle_left_transparency_texture[23][50] = 0;	doodle_left_transparency_texture[23][51] = 0;	doodle_left_transparency_texture[23][52] = 0;	doodle_left_transparency_texture[23][53] = 0;	doodle_left_transparency_texture[23][54] = 0;	doodle_left_transparency_texture[23][55] = 0;	doodle_left_transparency_texture[23][56] = 0;	doodle_left_transparency_texture[23][57] = 0;	doodle_left_transparency_texture[23][58] = 0;	doodle_left_transparency_texture[23][59] = 0;	doodle_left_transparency_texture[23][60] = 0;	doodle_left_transparency_texture[23][61] = 0;	doodle_left_transparency_texture[23][62] = 0;	doodle_left_transparency_texture[23][63] = 0;	doodle_left_transparency_texture[23][64] = 0;	doodle_left_transparency_texture[23][65] = 0;	doodle_left_transparency_texture[23][66] = 0;	doodle_left_transparency_texture[23][67] = 0;	doodle_left_transparency_texture[23][68] = 0;	doodle_left_transparency_texture[23][69] = 0;	doodle_left_transparency_texture[23][70] = 0;	doodle_left_transparency_texture[23][71] = 0;	doodle_left_transparency_texture[23][72] = 0;	doodle_left_transparency_texture[23][73] = 0;	doodle_left_transparency_texture[23][74] = 0;	doodle_left_transparency_texture[23][75] = 0;	doodle_left_transparency_texture[23][76] = 1;	doodle_left_transparency_texture[23][77] = 1;	doodle_left_transparency_texture[23][78] = 1;	doodle_left_transparency_texture[23][79] = 1;	doodle_left_transparency_texture[24][0] = 1;	doodle_left_transparency_texture[24][1] = 1;	doodle_left_transparency_texture[24][2] = 1;	doodle_left_transparency_texture[24][3] = 1;	doodle_left_transparency_texture[24][4] = 0;	doodle_left_transparency_texture[24][5] = 0;	doodle_left_transparency_texture[24][6] = 0;	doodle_left_transparency_texture[24][7] = 0;	doodle_left_transparency_texture[24][8] = 0;	doodle_left_transparency_texture[24][9] = 0;	doodle_left_transparency_texture[24][10] = 0;	doodle_left_transparency_texture[24][11] = 0;	doodle_left_transparency_texture[24][12] = 0;	doodle_left_transparency_texture[24][13] = 0;	doodle_left_transparency_texture[24][14] = 0;	doodle_left_transparency_texture[24][15] = 0;	doodle_left_transparency_texture[24][16] = 0;	doodle_left_transparency_texture[24][17] = 0;	doodle_left_transparency_texture[24][18] = 0;	doodle_left_transparency_texture[24][19] = 0;	doodle_left_transparency_texture[24][20] = 0;	doodle_left_transparency_texture[24][21] = 0;	doodle_left_transparency_texture[24][22] = 0;	doodle_left_transparency_texture[24][23] = 0;	doodle_left_transparency_texture[24][24] = 0;	doodle_left_transparency_texture[24][25] = 0;	doodle_left_transparency_texture[24][26] = 0;	doodle_left_transparency_texture[24][27] = 0;	doodle_left_transparency_texture[24][28] = 0;	doodle_left_transparency_texture[24][29] = 0;	doodle_left_transparency_texture[24][30] = 0;	doodle_left_transparency_texture[24][31] = 0;	doodle_left_transparency_texture[24][32] = 0;	doodle_left_transparency_texture[24][33] = 0;	doodle_left_transparency_texture[24][34] = 0;	doodle_left_transparency_texture[24][35] = 0;	doodle_left_transparency_texture[24][36] = 0;	doodle_left_transparency_texture[24][37] = 0;	doodle_left_transparency_texture[24][38] = 0;	doodle_left_transparency_texture[24][39] = 0;	doodle_left_transparency_texture[24][40] = 0;	doodle_left_transparency_texture[24][41] = 0;	doodle_left_transparency_texture[24][42] = 0;	doodle_left_transparency_texture[24][43] = 0;	doodle_left_transparency_texture[24][44] = 0;	doodle_left_transparency_texture[24][45] = 0;	doodle_left_transparency_texture[24][46] = 0;	doodle_left_transparency_texture[24][47] = 0;	doodle_left_transparency_texture[24][48] = 0;	doodle_left_transparency_texture[24][49] = 0;	doodle_left_transparency_texture[24][50] = 0;	doodle_left_transparency_texture[24][51] = 0;	doodle_left_transparency_texture[24][52] = 0;	doodle_left_transparency_texture[24][53] = 0;	doodle_left_transparency_texture[24][54] = 0;	doodle_left_transparency_texture[24][55] = 0;	doodle_left_transparency_texture[24][56] = 0;	doodle_left_transparency_texture[24][57] = 0;	doodle_left_transparency_texture[24][58] = 0;	doodle_left_transparency_texture[24][59] = 0;	doodle_left_transparency_texture[24][60] = 0;	doodle_left_transparency_texture[24][61] = 0;	doodle_left_transparency_texture[24][62] = 0;	doodle_left_transparency_texture[24][63] = 0;	doodle_left_transparency_texture[24][64] = 0;	doodle_left_transparency_texture[24][65] = 0;	doodle_left_transparency_texture[24][66] = 0;	doodle_left_transparency_texture[24][67] = 0;	doodle_left_transparency_texture[24][68] = 0;	doodle_left_transparency_texture[24][69] = 0;	doodle_left_transparency_texture[24][70] = 0;	doodle_left_transparency_texture[24][71] = 0;	doodle_left_transparency_texture[24][72] = 0;	doodle_left_transparency_texture[24][73] = 0;	doodle_left_transparency_texture[24][74] = 0;	doodle_left_transparency_texture[24][75] = 0;	doodle_left_transparency_texture[24][76] = 1;	doodle_left_transparency_texture[24][77] = 1;	doodle_left_transparency_texture[24][78] = 1;	doodle_left_transparency_texture[24][79] = 1;	doodle_left_transparency_texture[25][0] = 1;	doodle_left_transparency_texture[25][1] = 1;	doodle_left_transparency_texture[25][2] = 1;	doodle_left_transparency_texture[25][3] = 1;	doodle_left_transparency_texture[25][4] = 0;	doodle_left_transparency_texture[25][5] = 0;	doodle_left_transparency_texture[25][6] = 0;	doodle_left_transparency_texture[25][7] = 0;	doodle_left_transparency_texture[25][8] = 0;	doodle_left_transparency_texture[25][9] = 0;	doodle_left_transparency_texture[25][10] = 0;	doodle_left_transparency_texture[25][11] = 0;	doodle_left_transparency_texture[25][12] = 0;	doodle_left_transparency_texture[25][13] = 0;	doodle_left_transparency_texture[25][14] = 0;	doodle_left_transparency_texture[25][15] = 0;	doodle_left_transparency_texture[25][16] = 0;	doodle_left_transparency_texture[25][17] = 0;	doodle_left_transparency_texture[25][18] = 0;	doodle_left_transparency_texture[25][19] = 0;	doodle_left_transparency_texture[25][20] = 0;	doodle_left_transparency_texture[25][21] = 0;	doodle_left_transparency_texture[25][22] = 0;	doodle_left_transparency_texture[25][23] = 0;	doodle_left_transparency_texture[25][24] = 0;	doodle_left_transparency_texture[25][25] = 0;	doodle_left_transparency_texture[25][26] = 0;	doodle_left_transparency_texture[25][27] = 0;	doodle_left_transparency_texture[25][28] = 0;	doodle_left_transparency_texture[25][29] = 0;	doodle_left_transparency_texture[25][30] = 0;	doodle_left_transparency_texture[25][31] = 0;	doodle_left_transparency_texture[25][32] = 0;	doodle_left_transparency_texture[25][33] = 0;	doodle_left_transparency_texture[25][34] = 0;	doodle_left_transparency_texture[25][35] = 0;	doodle_left_transparency_texture[25][36] = 0;	doodle_left_transparency_texture[25][37] = 0;	doodle_left_transparency_texture[25][38] = 0;	doodle_left_transparency_texture[25][39] = 0;	doodle_left_transparency_texture[25][40] = 0;	doodle_left_transparency_texture[25][41] = 0;	doodle_left_transparency_texture[25][42] = 0;	doodle_left_transparency_texture[25][43] = 0;	doodle_left_transparency_texture[25][44] = 0;	doodle_left_transparency_texture[25][45] = 0;	doodle_left_transparency_texture[25][46] = 0;	doodle_left_transparency_texture[25][47] = 0;	doodle_left_transparency_texture[25][48] = 0;	doodle_left_transparency_texture[25][49] = 0;	doodle_left_transparency_texture[25][50] = 0;	doodle_left_transparency_texture[25][51] = 0;	doodle_left_transparency_texture[25][52] = 0;	doodle_left_transparency_texture[25][53] = 0;	doodle_left_transparency_texture[25][54] = 0;	doodle_left_transparency_texture[25][55] = 0;	doodle_left_transparency_texture[25][56] = 0;	doodle_left_transparency_texture[25][57] = 0;	doodle_left_transparency_texture[25][58] = 0;	doodle_left_transparency_texture[25][59] = 0;	doodle_left_transparency_texture[25][60] = 0;	doodle_left_transparency_texture[25][61] = 0;	doodle_left_transparency_texture[25][62] = 0;	doodle_left_transparency_texture[25][63] = 0;	doodle_left_transparency_texture[25][64] = 0;	doodle_left_transparency_texture[25][65] = 0;	doodle_left_transparency_texture[25][66] = 0;	doodle_left_transparency_texture[25][67] = 0;	doodle_left_transparency_texture[25][68] = 0;	doodle_left_transparency_texture[25][69] = 0;	doodle_left_transparency_texture[25][70] = 0;	doodle_left_transparency_texture[25][71] = 0;	doodle_left_transparency_texture[25][72] = 0;	doodle_left_transparency_texture[25][73] = 0;	doodle_left_transparency_texture[25][74] = 0;	doodle_left_transparency_texture[25][75] = 0;	doodle_left_transparency_texture[25][76] = 1;	doodle_left_transparency_texture[25][77] = 1;	doodle_left_transparency_texture[25][78] = 1;	doodle_left_transparency_texture[25][79] = 1;	doodle_left_transparency_texture[26][0] = 1;	doodle_left_transparency_texture[26][1] = 1;	doodle_left_transparency_texture[26][2] = 1;	doodle_left_transparency_texture[26][3] = 1;	doodle_left_transparency_texture[26][4] = 0;	doodle_left_transparency_texture[26][5] = 0;	doodle_left_transparency_texture[26][6] = 0;	doodle_left_transparency_texture[26][7] = 0;	doodle_left_transparency_texture[26][8] = 0;	doodle_left_transparency_texture[26][9] = 0;	doodle_left_transparency_texture[26][10] = 0;	doodle_left_transparency_texture[26][11] = 0;	doodle_left_transparency_texture[26][12] = 0;	doodle_left_transparency_texture[26][13] = 0;	doodle_left_transparency_texture[26][14] = 0;	doodle_left_transparency_texture[26][15] = 0;	doodle_left_transparency_texture[26][16] = 0;	doodle_left_transparency_texture[26][17] = 0;	doodle_left_transparency_texture[26][18] = 0;	doodle_left_transparency_texture[26][19] = 0;	doodle_left_transparency_texture[26][20] = 0;	doodle_left_transparency_texture[26][21] = 0;	doodle_left_transparency_texture[26][22] = 0;	doodle_left_transparency_texture[26][23] = 0;	doodle_left_transparency_texture[26][24] = 0;	doodle_left_transparency_texture[26][25] = 0;	doodle_left_transparency_texture[26][26] = 0;	doodle_left_transparency_texture[26][27] = 0;	doodle_left_transparency_texture[26][28] = 0;	doodle_left_transparency_texture[26][29] = 0;	doodle_left_transparency_texture[26][30] = 0;	doodle_left_transparency_texture[26][31] = 0;	doodle_left_transparency_texture[26][32] = 0;	doodle_left_transparency_texture[26][33] = 0;	doodle_left_transparency_texture[26][34] = 0;	doodle_left_transparency_texture[26][35] = 0;	doodle_left_transparency_texture[26][36] = 0;	doodle_left_transparency_texture[26][37] = 0;	doodle_left_transparency_texture[26][38] = 0;	doodle_left_transparency_texture[26][39] = 0;	doodle_left_transparency_texture[26][40] = 0;	doodle_left_transparency_texture[26][41] = 0;	doodle_left_transparency_texture[26][42] = 0;	doodle_left_transparency_texture[26][43] = 0;	doodle_left_transparency_texture[26][44] = 0;	doodle_left_transparency_texture[26][45] = 0;	doodle_left_transparency_texture[26][46] = 0;	doodle_left_transparency_texture[26][47] = 0;	doodle_left_transparency_texture[26][48] = 0;	doodle_left_transparency_texture[26][49] = 0;	doodle_left_transparency_texture[26][50] = 0;	doodle_left_transparency_texture[26][51] = 0;	doodle_left_transparency_texture[26][52] = 0;	doodle_left_transparency_texture[26][53] = 0;	doodle_left_transparency_texture[26][54] = 0;	doodle_left_transparency_texture[26][55] = 0;	doodle_left_transparency_texture[26][56] = 0;	doodle_left_transparency_texture[26][57] = 0;	doodle_left_transparency_texture[26][58] = 0;	doodle_left_transparency_texture[26][59] = 0;	doodle_left_transparency_texture[26][60] = 0;	doodle_left_transparency_texture[26][61] = 0;	doodle_left_transparency_texture[26][62] = 0;	doodle_left_transparency_texture[26][63] = 0;	doodle_left_transparency_texture[26][64] = 0;	doodle_left_transparency_texture[26][65] = 0;	doodle_left_transparency_texture[26][66] = 0;	doodle_left_transparency_texture[26][67] = 0;	doodle_left_transparency_texture[26][68] = 0;	doodle_left_transparency_texture[26][69] = 0;	doodle_left_transparency_texture[26][70] = 0;	doodle_left_transparency_texture[26][71] = 0;	doodle_left_transparency_texture[26][72] = 0;	doodle_left_transparency_texture[26][73] = 0;	doodle_left_transparency_texture[26][74] = 0;	doodle_left_transparency_texture[26][75] = 0;	doodle_left_transparency_texture[26][76] = 1;	doodle_left_transparency_texture[26][77] = 1;	doodle_left_transparency_texture[26][78] = 1;	doodle_left_transparency_texture[26][79] = 1;	doodle_left_transparency_texture[27][0] = 1;	doodle_left_transparency_texture[27][1] = 1;	doodle_left_transparency_texture[27][2] = 1;	doodle_left_transparency_texture[27][3] = 1;	doodle_left_transparency_texture[27][4] = 0;	doodle_left_transparency_texture[27][5] = 0;	doodle_left_transparency_texture[27][6] = 0;	doodle_left_transparency_texture[27][7] = 0;	doodle_left_transparency_texture[27][8] = 0;	doodle_left_transparency_texture[27][9] = 0;	doodle_left_transparency_texture[27][10] = 0;	doodle_left_transparency_texture[27][11] = 0;	doodle_left_transparency_texture[27][12] = 0;	doodle_left_transparency_texture[27][13] = 0;	doodle_left_transparency_texture[27][14] = 0;	doodle_left_transparency_texture[27][15] = 0;	doodle_left_transparency_texture[27][16] = 0;	doodle_left_transparency_texture[27][17] = 0;	doodle_left_transparency_texture[27][18] = 0;	doodle_left_transparency_texture[27][19] = 0;	doodle_left_transparency_texture[27][20] = 0;	doodle_left_transparency_texture[27][21] = 0;	doodle_left_transparency_texture[27][22] = 0;	doodle_left_transparency_texture[27][23] = 0;	doodle_left_transparency_texture[27][24] = 0;	doodle_left_transparency_texture[27][25] = 0;	doodle_left_transparency_texture[27][26] = 0;	doodle_left_transparency_texture[27][27] = 0;	doodle_left_transparency_texture[27][28] = 0;	doodle_left_transparency_texture[27][29] = 0;	doodle_left_transparency_texture[27][30] = 0;	doodle_left_transparency_texture[27][31] = 0;	doodle_left_transparency_texture[27][32] = 0;	doodle_left_transparency_texture[27][33] = 0;	doodle_left_transparency_texture[27][34] = 0;	doodle_left_transparency_texture[27][35] = 0;	doodle_left_transparency_texture[27][36] = 0;	doodle_left_transparency_texture[27][37] = 0;	doodle_left_transparency_texture[27][38] = 0;	doodle_left_transparency_texture[27][39] = 0;	doodle_left_transparency_texture[27][40] = 0;	doodle_left_transparency_texture[27][41] = 0;	doodle_left_transparency_texture[27][42] = 0;	doodle_left_transparency_texture[27][43] = 0;	doodle_left_transparency_texture[27][44] = 0;	doodle_left_transparency_texture[27][45] = 0;	doodle_left_transparency_texture[27][46] = 0;	doodle_left_transparency_texture[27][47] = 0;	doodle_left_transparency_texture[27][48] = 0;	doodle_left_transparency_texture[27][49] = 0;	doodle_left_transparency_texture[27][50] = 0;	doodle_left_transparency_texture[27][51] = 0;	doodle_left_transparency_texture[27][52] = 0;	doodle_left_transparency_texture[27][53] = 0;	doodle_left_transparency_texture[27][54] = 0;	doodle_left_transparency_texture[27][55] = 0;	doodle_left_transparency_texture[27][56] = 0;	doodle_left_transparency_texture[27][57] = 0;	doodle_left_transparency_texture[27][58] = 0;	doodle_left_transparency_texture[27][59] = 0;	doodle_left_transparency_texture[27][60] = 0;	doodle_left_transparency_texture[27][61] = 0;	doodle_left_transparency_texture[27][62] = 0;	doodle_left_transparency_texture[27][63] = 0;	doodle_left_transparency_texture[27][64] = 0;	doodle_left_transparency_texture[27][65] = 0;	doodle_left_transparency_texture[27][66] = 0;	doodle_left_transparency_texture[27][67] = 0;	doodle_left_transparency_texture[27][68] = 0;	doodle_left_transparency_texture[27][69] = 0;	doodle_left_transparency_texture[27][70] = 0;	doodle_left_transparency_texture[27][71] = 0;	doodle_left_transparency_texture[27][72] = 0;	doodle_left_transparency_texture[27][73] = 0;	doodle_left_transparency_texture[27][74] = 0;	doodle_left_transparency_texture[27][75] = 0;	doodle_left_transparency_texture[27][76] = 1;	doodle_left_transparency_texture[27][77] = 1;	doodle_left_transparency_texture[27][78] = 1;	doodle_left_transparency_texture[27][79] = 1;	doodle_left_transparency_texture[28][0] = 1;	doodle_left_transparency_texture[28][1] = 1;	doodle_left_transparency_texture[28][2] = 1;	doodle_left_transparency_texture[28][3] = 1;	doodle_left_transparency_texture[28][4] = 0;	doodle_left_transparency_texture[28][5] = 0;	doodle_left_transparency_texture[28][6] = 0;	doodle_left_transparency_texture[28][7] = 0;	doodle_left_transparency_texture[28][8] = 0;	doodle_left_transparency_texture[28][9] = 0;	doodle_left_transparency_texture[28][10] = 0;	doodle_left_transparency_texture[28][11] = 0;	doodle_left_transparency_texture[28][12] = 0;	doodle_left_transparency_texture[28][13] = 0;	doodle_left_transparency_texture[28][14] = 0;	doodle_left_transparency_texture[28][15] = 0;	doodle_left_transparency_texture[28][16] = 0;	doodle_left_transparency_texture[28][17] = 0;	doodle_left_transparency_texture[28][18] = 0;	doodle_left_transparency_texture[28][19] = 0;	doodle_left_transparency_texture[28][20] = 0;	doodle_left_transparency_texture[28][21] = 0;	doodle_left_transparency_texture[28][22] = 0;	doodle_left_transparency_texture[28][23] = 0;	doodle_left_transparency_texture[28][24] = 0;	doodle_left_transparency_texture[28][25] = 0;	doodle_left_transparency_texture[28][26] = 0;	doodle_left_transparency_texture[28][27] = 0;	doodle_left_transparency_texture[28][28] = 0;	doodle_left_transparency_texture[28][29] = 0;	doodle_left_transparency_texture[28][30] = 0;	doodle_left_transparency_texture[28][31] = 0;	doodle_left_transparency_texture[28][32] = 0;	doodle_left_transparency_texture[28][33] = 0;	doodle_left_transparency_texture[28][34] = 0;	doodle_left_transparency_texture[28][35] = 0;	doodle_left_transparency_texture[28][36] = 0;	doodle_left_transparency_texture[28][37] = 0;	doodle_left_transparency_texture[28][38] = 0;	doodle_left_transparency_texture[28][39] = 0;	doodle_left_transparency_texture[28][40] = 0;	doodle_left_transparency_texture[28][41] = 0;	doodle_left_transparency_texture[28][42] = 0;	doodle_left_transparency_texture[28][43] = 0;	doodle_left_transparency_texture[28][44] = 0;	doodle_left_transparency_texture[28][45] = 0;	doodle_left_transparency_texture[28][46] = 0;	doodle_left_transparency_texture[28][47] = 0;	doodle_left_transparency_texture[28][48] = 0;	doodle_left_transparency_texture[28][49] = 0;	doodle_left_transparency_texture[28][50] = 0;	doodle_left_transparency_texture[28][51] = 0;	doodle_left_transparency_texture[28][52] = 0;	doodle_left_transparency_texture[28][53] = 0;	doodle_left_transparency_texture[28][54] = 0;	doodle_left_transparency_texture[28][55] = 0;	doodle_left_transparency_texture[28][56] = 0;	doodle_left_transparency_texture[28][57] = 0;	doodle_left_transparency_texture[28][58] = 0;	doodle_left_transparency_texture[28][59] = 0;	doodle_left_transparency_texture[28][60] = 0;	doodle_left_transparency_texture[28][61] = 0;	doodle_left_transparency_texture[28][62] = 0;	doodle_left_transparency_texture[28][63] = 0;	doodle_left_transparency_texture[28][64] = 0;	doodle_left_transparency_texture[28][65] = 0;	doodle_left_transparency_texture[28][66] = 0;	doodle_left_transparency_texture[28][67] = 0;	doodle_left_transparency_texture[28][68] = 0;	doodle_left_transparency_texture[28][69] = 0;	doodle_left_transparency_texture[28][70] = 0;	doodle_left_transparency_texture[28][71] = 0;	doodle_left_transparency_texture[28][72] = 0;	doodle_left_transparency_texture[28][73] = 0;	doodle_left_transparency_texture[28][74] = 0;	doodle_left_transparency_texture[28][75] = 0;	doodle_left_transparency_texture[28][76] = 1;	doodle_left_transparency_texture[28][77] = 1;	doodle_left_transparency_texture[28][78] = 1;	doodle_left_transparency_texture[28][79] = 1;	doodle_left_transparency_texture[29][0] = 1;	doodle_left_transparency_texture[29][1] = 1;	doodle_left_transparency_texture[29][2] = 1;	doodle_left_transparency_texture[29][3] = 1;	doodle_left_transparency_texture[29][4] = 0;	doodle_left_transparency_texture[29][5] = 0;	doodle_left_transparency_texture[29][6] = 0;	doodle_left_transparency_texture[29][7] = 0;	doodle_left_transparency_texture[29][8] = 0;	doodle_left_transparency_texture[29][9] = 0;	doodle_left_transparency_texture[29][10] = 0;	doodle_left_transparency_texture[29][11] = 0;	doodle_left_transparency_texture[29][12] = 0;	doodle_left_transparency_texture[29][13] = 0;	doodle_left_transparency_texture[29][14] = 0;	doodle_left_transparency_texture[29][15] = 0;	doodle_left_transparency_texture[29][16] = 0;	doodle_left_transparency_texture[29][17] = 0;	doodle_left_transparency_texture[29][18] = 0;	doodle_left_transparency_texture[29][19] = 0;	doodle_left_transparency_texture[29][20] = 0;	doodle_left_transparency_texture[29][21] = 0;	doodle_left_transparency_texture[29][22] = 0;	doodle_left_transparency_texture[29][23] = 0;	doodle_left_transparency_texture[29][24] = 0;	doodle_left_transparency_texture[29][25] = 0;	doodle_left_transparency_texture[29][26] = 0;	doodle_left_transparency_texture[29][27] = 0;	doodle_left_transparency_texture[29][28] = 0;	doodle_left_transparency_texture[29][29] = 0;	doodle_left_transparency_texture[29][30] = 0;	doodle_left_transparency_texture[29][31] = 0;	doodle_left_transparency_texture[29][32] = 0;	doodle_left_transparency_texture[29][33] = 0;	doodle_left_transparency_texture[29][34] = 0;	doodle_left_transparency_texture[29][35] = 0;	doodle_left_transparency_texture[29][36] = 0;	doodle_left_transparency_texture[29][37] = 0;	doodle_left_transparency_texture[29][38] = 0;	doodle_left_transparency_texture[29][39] = 0;	doodle_left_transparency_texture[29][40] = 0;	doodle_left_transparency_texture[29][41] = 0;	doodle_left_transparency_texture[29][42] = 0;	doodle_left_transparency_texture[29][43] = 0;	doodle_left_transparency_texture[29][44] = 0;	doodle_left_transparency_texture[29][45] = 0;	doodle_left_transparency_texture[29][46] = 0;	doodle_left_transparency_texture[29][47] = 0;	doodle_left_transparency_texture[29][48] = 0;	doodle_left_transparency_texture[29][49] = 0;	doodle_left_transparency_texture[29][50] = 0;	doodle_left_transparency_texture[29][51] = 0;	doodle_left_transparency_texture[29][52] = 0;	doodle_left_transparency_texture[29][53] = 0;	doodle_left_transparency_texture[29][54] = 0;	doodle_left_transparency_texture[29][55] = 0;	doodle_left_transparency_texture[29][56] = 0;	doodle_left_transparency_texture[29][57] = 0;	doodle_left_transparency_texture[29][58] = 0;	doodle_left_transparency_texture[29][59] = 0;	doodle_left_transparency_texture[29][60] = 0;	doodle_left_transparency_texture[29][61] = 0;	doodle_left_transparency_texture[29][62] = 0;	doodle_left_transparency_texture[29][63] = 0;	doodle_left_transparency_texture[29][64] = 0;	doodle_left_transparency_texture[29][65] = 0;	doodle_left_transparency_texture[29][66] = 0;	doodle_left_transparency_texture[29][67] = 0;	doodle_left_transparency_texture[29][68] = 0;	doodle_left_transparency_texture[29][69] = 0;	doodle_left_transparency_texture[29][70] = 0;	doodle_left_transparency_texture[29][71] = 0;	doodle_left_transparency_texture[29][72] = 0;	doodle_left_transparency_texture[29][73] = 0;	doodle_left_transparency_texture[29][74] = 0;	doodle_left_transparency_texture[29][75] = 0;	doodle_left_transparency_texture[29][76] = 1;	doodle_left_transparency_texture[29][77] = 1;	doodle_left_transparency_texture[29][78] = 1;	doodle_left_transparency_texture[29][79] = 1;	doodle_left_transparency_texture[30][0] = 1;	doodle_left_transparency_texture[30][1] = 1;	doodle_left_transparency_texture[30][2] = 1;	doodle_left_transparency_texture[30][3] = 1;	doodle_left_transparency_texture[30][4] = 0;	doodle_left_transparency_texture[30][5] = 0;	doodle_left_transparency_texture[30][6] = 0;	doodle_left_transparency_texture[30][7] = 0;	doodle_left_transparency_texture[30][8] = 0;	doodle_left_transparency_texture[30][9] = 0;	doodle_left_transparency_texture[30][10] = 0;	doodle_left_transparency_texture[30][11] = 0;	doodle_left_transparency_texture[30][12] = 0;	doodle_left_transparency_texture[30][13] = 0;	doodle_left_transparency_texture[30][14] = 0;	doodle_left_transparency_texture[30][15] = 0;	doodle_left_transparency_texture[30][16] = 0;	doodle_left_transparency_texture[30][17] = 0;	doodle_left_transparency_texture[30][18] = 0;	doodle_left_transparency_texture[30][19] = 0;	doodle_left_transparency_texture[30][20] = 0;	doodle_left_transparency_texture[30][21] = 0;	doodle_left_transparency_texture[30][22] = 0;	doodle_left_transparency_texture[30][23] = 0;	doodle_left_transparency_texture[30][24] = 0;	doodle_left_transparency_texture[30][25] = 0;	doodle_left_transparency_texture[30][26] = 0;	doodle_left_transparency_texture[30][27] = 0;	doodle_left_transparency_texture[30][28] = 0;	doodle_left_transparency_texture[30][29] = 0;	doodle_left_transparency_texture[30][30] = 0;	doodle_left_transparency_texture[30][31] = 0;	doodle_left_transparency_texture[30][32] = 0;	doodle_left_transparency_texture[30][33] = 0;	doodle_left_transparency_texture[30][34] = 0;	doodle_left_transparency_texture[30][35] = 0;	doodle_left_transparency_texture[30][36] = 0;	doodle_left_transparency_texture[30][37] = 0;	doodle_left_transparency_texture[30][38] = 0;	doodle_left_transparency_texture[30][39] = 0;	doodle_left_transparency_texture[30][40] = 0;	doodle_left_transparency_texture[30][41] = 0;	doodle_left_transparency_texture[30][42] = 0;	doodle_left_transparency_texture[30][43] = 0;	doodle_left_transparency_texture[30][44] = 0;	doodle_left_transparency_texture[30][45] = 0;	doodle_left_transparency_texture[30][46] = 0;	doodle_left_transparency_texture[30][47] = 0;	doodle_left_transparency_texture[30][48] = 0;	doodle_left_transparency_texture[30][49] = 0;	doodle_left_transparency_texture[30][50] = 0;	doodle_left_transparency_texture[30][51] = 0;	doodle_left_transparency_texture[30][52] = 0;	doodle_left_transparency_texture[30][53] = 0;	doodle_left_transparency_texture[30][54] = 0;	doodle_left_transparency_texture[30][55] = 0;	doodle_left_transparency_texture[30][56] = 0;	doodle_left_transparency_texture[30][57] = 0;	doodle_left_transparency_texture[30][58] = 0;	doodle_left_transparency_texture[30][59] = 0;	doodle_left_transparency_texture[30][60] = 0;	doodle_left_transparency_texture[30][61] = 0;	doodle_left_transparency_texture[30][62] = 0;	doodle_left_transparency_texture[30][63] = 0;	doodle_left_transparency_texture[30][64] = 0;	doodle_left_transparency_texture[30][65] = 0;	doodle_left_transparency_texture[30][66] = 0;	doodle_left_transparency_texture[30][67] = 0;	doodle_left_transparency_texture[30][68] = 0;	doodle_left_transparency_texture[30][69] = 0;	doodle_left_transparency_texture[30][70] = 0;	doodle_left_transparency_texture[30][71] = 0;	doodle_left_transparency_texture[30][72] = 0;	doodle_left_transparency_texture[30][73] = 0;	doodle_left_transparency_texture[30][74] = 0;	doodle_left_transparency_texture[30][75] = 0;	doodle_left_transparency_texture[30][76] = 1;	doodle_left_transparency_texture[30][77] = 1;	doodle_left_transparency_texture[30][78] = 1;	doodle_left_transparency_texture[30][79] = 1;	doodle_left_transparency_texture[31][0] = 1;	doodle_left_transparency_texture[31][1] = 1;	doodle_left_transparency_texture[31][2] = 1;	doodle_left_transparency_texture[31][3] = 1;	doodle_left_transparency_texture[31][4] = 0;	doodle_left_transparency_texture[31][5] = 0;	doodle_left_transparency_texture[31][6] = 0;	doodle_left_transparency_texture[31][7] = 0;	doodle_left_transparency_texture[31][8] = 0;	doodle_left_transparency_texture[31][9] = 0;	doodle_left_transparency_texture[31][10] = 0;	doodle_left_transparency_texture[31][11] = 0;	doodle_left_transparency_texture[31][12] = 0;	doodle_left_transparency_texture[31][13] = 0;	doodle_left_transparency_texture[31][14] = 0;	doodle_left_transparency_texture[31][15] = 0;	doodle_left_transparency_texture[31][16] = 0;	doodle_left_transparency_texture[31][17] = 0;	doodle_left_transparency_texture[31][18] = 0;	doodle_left_transparency_texture[31][19] = 0;	doodle_left_transparency_texture[31][20] = 0;	doodle_left_transparency_texture[31][21] = 0;	doodle_left_transparency_texture[31][22] = 0;	doodle_left_transparency_texture[31][23] = 0;	doodle_left_transparency_texture[31][24] = 0;	doodle_left_transparency_texture[31][25] = 0;	doodle_left_transparency_texture[31][26] = 0;	doodle_left_transparency_texture[31][27] = 0;	doodle_left_transparency_texture[31][28] = 0;	doodle_left_transparency_texture[31][29] = 0;	doodle_left_transparency_texture[31][30] = 0;	doodle_left_transparency_texture[31][31] = 0;	doodle_left_transparency_texture[31][32] = 0;	doodle_left_transparency_texture[31][33] = 0;	doodle_left_transparency_texture[31][34] = 0;	doodle_left_transparency_texture[31][35] = 0;	doodle_left_transparency_texture[31][36] = 0;	doodle_left_transparency_texture[31][37] = 0;	doodle_left_transparency_texture[31][38] = 0;	doodle_left_transparency_texture[31][39] = 0;	doodle_left_transparency_texture[31][40] = 0;	doodle_left_transparency_texture[31][41] = 0;	doodle_left_transparency_texture[31][42] = 0;	doodle_left_transparency_texture[31][43] = 0;	doodle_left_transparency_texture[31][44] = 0;	doodle_left_transparency_texture[31][45] = 0;	doodle_left_transparency_texture[31][46] = 0;	doodle_left_transparency_texture[31][47] = 0;	doodle_left_transparency_texture[31][48] = 0;	doodle_left_transparency_texture[31][49] = 0;	doodle_left_transparency_texture[31][50] = 0;	doodle_left_transparency_texture[31][51] = 0;	doodle_left_transparency_texture[31][52] = 0;	doodle_left_transparency_texture[31][53] = 0;	doodle_left_transparency_texture[31][54] = 0;	doodle_left_transparency_texture[31][55] = 0;	doodle_left_transparency_texture[31][56] = 0;	doodle_left_transparency_texture[31][57] = 0;	doodle_left_transparency_texture[31][58] = 0;	doodle_left_transparency_texture[31][59] = 0;	doodle_left_transparency_texture[31][60] = 0;	doodle_left_transparency_texture[31][61] = 0;	doodle_left_transparency_texture[31][62] = 0;	doodle_left_transparency_texture[31][63] = 0;	doodle_left_transparency_texture[31][64] = 0;	doodle_left_transparency_texture[31][65] = 0;	doodle_left_transparency_texture[31][66] = 0;	doodle_left_transparency_texture[31][67] = 0;	doodle_left_transparency_texture[31][68] = 0;	doodle_left_transparency_texture[31][69] = 0;	doodle_left_transparency_texture[31][70] = 0;	doodle_left_transparency_texture[31][71] = 0;	doodle_left_transparency_texture[31][72] = 0;	doodle_left_transparency_texture[31][73] = 0;	doodle_left_transparency_texture[31][74] = 0;	doodle_left_transparency_texture[31][75] = 0;	doodle_left_transparency_texture[31][76] = 1;	doodle_left_transparency_texture[31][77] = 1;	doodle_left_transparency_texture[31][78] = 1;	doodle_left_transparency_texture[31][79] = 1;	doodle_left_transparency_texture[32][0] = 1;	doodle_left_transparency_texture[32][1] = 1;	doodle_left_transparency_texture[32][2] = 1;	doodle_left_transparency_texture[32][3] = 1;	doodle_left_transparency_texture[32][4] = 0;	doodle_left_transparency_texture[32][5] = 0;	doodle_left_transparency_texture[32][6] = 0;	doodle_left_transparency_texture[32][7] = 0;	doodle_left_transparency_texture[32][8] = 0;	doodle_left_transparency_texture[32][9] = 0;	doodle_left_transparency_texture[32][10] = 0;	doodle_left_transparency_texture[32][11] = 0;	doodle_left_transparency_texture[32][12] = 0;	doodle_left_transparency_texture[32][13] = 0;	doodle_left_transparency_texture[32][14] = 0;	doodle_left_transparency_texture[32][15] = 0;	doodle_left_transparency_texture[32][16] = 0;	doodle_left_transparency_texture[32][17] = 0;	doodle_left_transparency_texture[32][18] = 0;	doodle_left_transparency_texture[32][19] = 0;	doodle_left_transparency_texture[32][20] = 0;	doodle_left_transparency_texture[32][21] = 0;	doodle_left_transparency_texture[32][22] = 0;	doodle_left_transparency_texture[32][23] = 0;	doodle_left_transparency_texture[32][24] = 0;	doodle_left_transparency_texture[32][25] = 0;	doodle_left_transparency_texture[32][26] = 0;	doodle_left_transparency_texture[32][27] = 0;	doodle_left_transparency_texture[32][28] = 0;	doodle_left_transparency_texture[32][29] = 0;	doodle_left_transparency_texture[32][30] = 0;	doodle_left_transparency_texture[32][31] = 0;	doodle_left_transparency_texture[32][32] = 0;	doodle_left_transparency_texture[32][33] = 0;	doodle_left_transparency_texture[32][34] = 0;	doodle_left_transparency_texture[32][35] = 0;	doodle_left_transparency_texture[32][36] = 0;	doodle_left_transparency_texture[32][37] = 0;	doodle_left_transparency_texture[32][38] = 0;	doodle_left_transparency_texture[32][39] = 0;	doodle_left_transparency_texture[32][40] = 0;	doodle_left_transparency_texture[32][41] = 0;	doodle_left_transparency_texture[32][42] = 0;	doodle_left_transparency_texture[32][43] = 0;	doodle_left_transparency_texture[32][44] = 0;	doodle_left_transparency_texture[32][45] = 0;	doodle_left_transparency_texture[32][46] = 0;	doodle_left_transparency_texture[32][47] = 0;	doodle_left_transparency_texture[32][48] = 0;	doodle_left_transparency_texture[32][49] = 0;	doodle_left_transparency_texture[32][50] = 0;	doodle_left_transparency_texture[32][51] = 0;	doodle_left_transparency_texture[32][52] = 0;	doodle_left_transparency_texture[32][53] = 0;	doodle_left_transparency_texture[32][54] = 0;	doodle_left_transparency_texture[32][55] = 0;	doodle_left_transparency_texture[32][56] = 0;	doodle_left_transparency_texture[32][57] = 0;	doodle_left_transparency_texture[32][58] = 0;	doodle_left_transparency_texture[32][59] = 0;	doodle_left_transparency_texture[32][60] = 0;	doodle_left_transparency_texture[32][61] = 0;	doodle_left_transparency_texture[32][62] = 0;	doodle_left_transparency_texture[32][63] = 0;	doodle_left_transparency_texture[32][64] = 0;	doodle_left_transparency_texture[32][65] = 0;	doodle_left_transparency_texture[32][66] = 0;	doodle_left_transparency_texture[32][67] = 0;	doodle_left_transparency_texture[32][68] = 0;	doodle_left_transparency_texture[32][69] = 0;	doodle_left_transparency_texture[32][70] = 0;	doodle_left_transparency_texture[32][71] = 0;	doodle_left_transparency_texture[32][72] = 0;	doodle_left_transparency_texture[32][73] = 0;	doodle_left_transparency_texture[32][74] = 0;	doodle_left_transparency_texture[32][75] = 0;	doodle_left_transparency_texture[32][76] = 1;	doodle_left_transparency_texture[32][77] = 1;	doodle_left_transparency_texture[32][78] = 1;	doodle_left_transparency_texture[32][79] = 1;	doodle_left_transparency_texture[33][0] = 1;	doodle_left_transparency_texture[33][1] = 1;	doodle_left_transparency_texture[33][2] = 1;	doodle_left_transparency_texture[33][3] = 1;	doodle_left_transparency_texture[33][4] = 0;	doodle_left_transparency_texture[33][5] = 0;	doodle_left_transparency_texture[33][6] = 0;	doodle_left_transparency_texture[33][7] = 0;	doodle_left_transparency_texture[33][8] = 0;	doodle_left_transparency_texture[33][9] = 0;	doodle_left_transparency_texture[33][10] = 0;	doodle_left_transparency_texture[33][11] = 0;	doodle_left_transparency_texture[33][12] = 0;	doodle_left_transparency_texture[33][13] = 0;	doodle_left_transparency_texture[33][14] = 0;	doodle_left_transparency_texture[33][15] = 0;	doodle_left_transparency_texture[33][16] = 0;	doodle_left_transparency_texture[33][17] = 0;	doodle_left_transparency_texture[33][18] = 0;	doodle_left_transparency_texture[33][19] = 0;	doodle_left_transparency_texture[33][20] = 0;	doodle_left_transparency_texture[33][21] = 0;	doodle_left_transparency_texture[33][22] = 0;	doodle_left_transparency_texture[33][23] = 0;	doodle_left_transparency_texture[33][24] = 0;	doodle_left_transparency_texture[33][25] = 0;	doodle_left_transparency_texture[33][26] = 0;	doodle_left_transparency_texture[33][27] = 0;	doodle_left_transparency_texture[33][28] = 0;	doodle_left_transparency_texture[33][29] = 0;	doodle_left_transparency_texture[33][30] = 0;	doodle_left_transparency_texture[33][31] = 0;	doodle_left_transparency_texture[33][32] = 0;	doodle_left_transparency_texture[33][33] = 0;	doodle_left_transparency_texture[33][34] = 0;	doodle_left_transparency_texture[33][35] = 0;	doodle_left_transparency_texture[33][36] = 0;	doodle_left_transparency_texture[33][37] = 0;	doodle_left_transparency_texture[33][38] = 0;	doodle_left_transparency_texture[33][39] = 0;	doodle_left_transparency_texture[33][40] = 0;	doodle_left_transparency_texture[33][41] = 0;	doodle_left_transparency_texture[33][42] = 0;	doodle_left_transparency_texture[33][43] = 0;	doodle_left_transparency_texture[33][44] = 0;	doodle_left_transparency_texture[33][45] = 0;	doodle_left_transparency_texture[33][46] = 0;	doodle_left_transparency_texture[33][47] = 0;	doodle_left_transparency_texture[33][48] = 0;	doodle_left_transparency_texture[33][49] = 0;	doodle_left_transparency_texture[33][50] = 0;	doodle_left_transparency_texture[33][51] = 0;	doodle_left_transparency_texture[33][52] = 0;	doodle_left_transparency_texture[33][53] = 0;	doodle_left_transparency_texture[33][54] = 0;	doodle_left_transparency_texture[33][55] = 0;	doodle_left_transparency_texture[33][56] = 0;	doodle_left_transparency_texture[33][57] = 0;	doodle_left_transparency_texture[33][58] = 0;	doodle_left_transparency_texture[33][59] = 0;	doodle_left_transparency_texture[33][60] = 0;	doodle_left_transparency_texture[33][61] = 0;	doodle_left_transparency_texture[33][62] = 0;	doodle_left_transparency_texture[33][63] = 0;	doodle_left_transparency_texture[33][64] = 0;	doodle_left_transparency_texture[33][65] = 0;	doodle_left_transparency_texture[33][66] = 0;	doodle_left_transparency_texture[33][67] = 0;	doodle_left_transparency_texture[33][68] = 0;	doodle_left_transparency_texture[33][69] = 0;	doodle_left_transparency_texture[33][70] = 0;	doodle_left_transparency_texture[33][71] = 0;	doodle_left_transparency_texture[33][72] = 0;	doodle_left_transparency_texture[33][73] = 0;	doodle_left_transparency_texture[33][74] = 0;	doodle_left_transparency_texture[33][75] = 0;	doodle_left_transparency_texture[33][76] = 1;	doodle_left_transparency_texture[33][77] = 1;	doodle_left_transparency_texture[33][78] = 1;	doodle_left_transparency_texture[33][79] = 1;	doodle_left_transparency_texture[34][0] = 1;	doodle_left_transparency_texture[34][1] = 1;	doodle_left_transparency_texture[34][2] = 1;	doodle_left_transparency_texture[34][3] = 1;	doodle_left_transparency_texture[34][4] = 0;	doodle_left_transparency_texture[34][5] = 0;	doodle_left_transparency_texture[34][6] = 0;	doodle_left_transparency_texture[34][7] = 0;	doodle_left_transparency_texture[34][8] = 0;	doodle_left_transparency_texture[34][9] = 0;	doodle_left_transparency_texture[34][10] = 0;	doodle_left_transparency_texture[34][11] = 0;	doodle_left_transparency_texture[34][12] = 0;	doodle_left_transparency_texture[34][13] = 0;	doodle_left_transparency_texture[34][14] = 0;	doodle_left_transparency_texture[34][15] = 0;	doodle_left_transparency_texture[34][16] = 0;	doodle_left_transparency_texture[34][17] = 0;	doodle_left_transparency_texture[34][18] = 0;	doodle_left_transparency_texture[34][19] = 0;	doodle_left_transparency_texture[34][20] = 0;	doodle_left_transparency_texture[34][21] = 0;	doodle_left_transparency_texture[34][22] = 0;	doodle_left_transparency_texture[34][23] = 0;	doodle_left_transparency_texture[34][24] = 0;	doodle_left_transparency_texture[34][25] = 0;	doodle_left_transparency_texture[34][26] = 0;	doodle_left_transparency_texture[34][27] = 0;	doodle_left_transparency_texture[34][28] = 0;	doodle_left_transparency_texture[34][29] = 0;	doodle_left_transparency_texture[34][30] = 0;	doodle_left_transparency_texture[34][31] = 0;	doodle_left_transparency_texture[34][32] = 0;	doodle_left_transparency_texture[34][33] = 0;	doodle_left_transparency_texture[34][34] = 0;	doodle_left_transparency_texture[34][35] = 0;	doodle_left_transparency_texture[34][36] = 0;	doodle_left_transparency_texture[34][37] = 0;	doodle_left_transparency_texture[34][38] = 0;	doodle_left_transparency_texture[34][39] = 0;	doodle_left_transparency_texture[34][40] = 0;	doodle_left_transparency_texture[34][41] = 0;	doodle_left_transparency_texture[34][42] = 0;	doodle_left_transparency_texture[34][43] = 0;	doodle_left_transparency_texture[34][44] = 0;	doodle_left_transparency_texture[34][45] = 0;	doodle_left_transparency_texture[34][46] = 0;	doodle_left_transparency_texture[34][47] = 0;	doodle_left_transparency_texture[34][48] = 0;	doodle_left_transparency_texture[34][49] = 0;	doodle_left_transparency_texture[34][50] = 0;	doodle_left_transparency_texture[34][51] = 0;	doodle_left_transparency_texture[34][52] = 0;	doodle_left_transparency_texture[34][53] = 0;	doodle_left_transparency_texture[34][54] = 0;	doodle_left_transparency_texture[34][55] = 0;	doodle_left_transparency_texture[34][56] = 0;	doodle_left_transparency_texture[34][57] = 0;	doodle_left_transparency_texture[34][58] = 0;	doodle_left_transparency_texture[34][59] = 0;	doodle_left_transparency_texture[34][60] = 0;	doodle_left_transparency_texture[34][61] = 0;	doodle_left_transparency_texture[34][62] = 0;	doodle_left_transparency_texture[34][63] = 0;	doodle_left_transparency_texture[34][64] = 0;	doodle_left_transparency_texture[34][65] = 0;	doodle_left_transparency_texture[34][66] = 0;	doodle_left_transparency_texture[34][67] = 0;	doodle_left_transparency_texture[34][68] = 0;	doodle_left_transparency_texture[34][69] = 0;	doodle_left_transparency_texture[34][70] = 0;	doodle_left_transparency_texture[34][71] = 0;	doodle_left_transparency_texture[34][72] = 0;	doodle_left_transparency_texture[34][73] = 0;	doodle_left_transparency_texture[34][74] = 0;	doodle_left_transparency_texture[34][75] = 0;	doodle_left_transparency_texture[34][76] = 1;	doodle_left_transparency_texture[34][77] = 1;	doodle_left_transparency_texture[34][78] = 1;	doodle_left_transparency_texture[34][79] = 1;	doodle_left_transparency_texture[35][0] = 1;	doodle_left_transparency_texture[35][1] = 1;	doodle_left_transparency_texture[35][2] = 1;	doodle_left_transparency_texture[35][3] = 1;	doodle_left_transparency_texture[35][4] = 0;	doodle_left_transparency_texture[35][5] = 0;	doodle_left_transparency_texture[35][6] = 0;	doodle_left_transparency_texture[35][7] = 0;	doodle_left_transparency_texture[35][8] = 0;	doodle_left_transparency_texture[35][9] = 0;	doodle_left_transparency_texture[35][10] = 0;	doodle_left_transparency_texture[35][11] = 0;	doodle_left_transparency_texture[35][12] = 0;	doodle_left_transparency_texture[35][13] = 0;	doodle_left_transparency_texture[35][14] = 0;	doodle_left_transparency_texture[35][15] = 0;	doodle_left_transparency_texture[35][16] = 0;	doodle_left_transparency_texture[35][17] = 0;	doodle_left_transparency_texture[35][18] = 0;	doodle_left_transparency_texture[35][19] = 0;	doodle_left_transparency_texture[35][20] = 0;	doodle_left_transparency_texture[35][21] = 0;	doodle_left_transparency_texture[35][22] = 0;	doodle_left_transparency_texture[35][23] = 0;	doodle_left_transparency_texture[35][24] = 0;	doodle_left_transparency_texture[35][25] = 0;	doodle_left_transparency_texture[35][26] = 0;	doodle_left_transparency_texture[35][27] = 0;	doodle_left_transparency_texture[35][28] = 0;	doodle_left_transparency_texture[35][29] = 0;	doodle_left_transparency_texture[35][30] = 0;	doodle_left_transparency_texture[35][31] = 0;	doodle_left_transparency_texture[35][32] = 0;	doodle_left_transparency_texture[35][33] = 0;	doodle_left_transparency_texture[35][34] = 0;	doodle_left_transparency_texture[35][35] = 0;	doodle_left_transparency_texture[35][36] = 0;	doodle_left_transparency_texture[35][37] = 0;	doodle_left_transparency_texture[35][38] = 0;	doodle_left_transparency_texture[35][39] = 0;	doodle_left_transparency_texture[35][40] = 0;	doodle_left_transparency_texture[35][41] = 0;	doodle_left_transparency_texture[35][42] = 0;	doodle_left_transparency_texture[35][43] = 0;	doodle_left_transparency_texture[35][44] = 0;	doodle_left_transparency_texture[35][45] = 0;	doodle_left_transparency_texture[35][46] = 0;	doodle_left_transparency_texture[35][47] = 0;	doodle_left_transparency_texture[35][48] = 0;	doodle_left_transparency_texture[35][49] = 0;	doodle_left_transparency_texture[35][50] = 0;	doodle_left_transparency_texture[35][51] = 0;	doodle_left_transparency_texture[35][52] = 0;	doodle_left_transparency_texture[35][53] = 0;	doodle_left_transparency_texture[35][54] = 0;	doodle_left_transparency_texture[35][55] = 0;	doodle_left_transparency_texture[35][56] = 0;	doodle_left_transparency_texture[35][57] = 0;	doodle_left_transparency_texture[35][58] = 0;	doodle_left_transparency_texture[35][59] = 0;	doodle_left_transparency_texture[35][60] = 0;	doodle_left_transparency_texture[35][61] = 0;	doodle_left_transparency_texture[35][62] = 0;	doodle_left_transparency_texture[35][63] = 0;	doodle_left_transparency_texture[35][64] = 0;	doodle_left_transparency_texture[35][65] = 0;	doodle_left_transparency_texture[35][66] = 0;	doodle_left_transparency_texture[35][67] = 0;	doodle_left_transparency_texture[35][68] = 0;	doodle_left_transparency_texture[35][69] = 0;	doodle_left_transparency_texture[35][70] = 0;	doodle_left_transparency_texture[35][71] = 0;	doodle_left_transparency_texture[35][72] = 0;	doodle_left_transparency_texture[35][73] = 0;	doodle_left_transparency_texture[35][74] = 0;	doodle_left_transparency_texture[35][75] = 0;	doodle_left_transparency_texture[35][76] = 1;	doodle_left_transparency_texture[35][77] = 1;	doodle_left_transparency_texture[35][78] = 1;	doodle_left_transparency_texture[35][79] = 1;	doodle_left_transparency_texture[36][0] = 1;	doodle_left_transparency_texture[36][1] = 1;	doodle_left_transparency_texture[36][2] = 1;	doodle_left_transparency_texture[36][3] = 1;	doodle_left_transparency_texture[36][4] = 1;	doodle_left_transparency_texture[36][5] = 1;	doodle_left_transparency_texture[36][6] = 1;	doodle_left_transparency_texture[36][7] = 1;	doodle_left_transparency_texture[36][8] = 1;	doodle_left_transparency_texture[36][9] = 1;	doodle_left_transparency_texture[36][10] = 1;	doodle_left_transparency_texture[36][11] = 1;	doodle_left_transparency_texture[36][12] = 1;	doodle_left_transparency_texture[36][13] = 1;	doodle_left_transparency_texture[36][14] = 1;	doodle_left_transparency_texture[36][15] = 1;	doodle_left_transparency_texture[36][16] = 1;	doodle_left_transparency_texture[36][17] = 1;	doodle_left_transparency_texture[36][18] = 1;	doodle_left_transparency_texture[36][19] = 1;	doodle_left_transparency_texture[36][20] = 1;	doodle_left_transparency_texture[36][21] = 1;	doodle_left_transparency_texture[36][22] = 1;	doodle_left_transparency_texture[36][23] = 1;	doodle_left_transparency_texture[36][24] = 1;	doodle_left_transparency_texture[36][25] = 1;	doodle_left_transparency_texture[36][26] = 1;	doodle_left_transparency_texture[36][27] = 1;	doodle_left_transparency_texture[36][28] = 0;	doodle_left_transparency_texture[36][29] = 0;	doodle_left_transparency_texture[36][30] = 0;	doodle_left_transparency_texture[36][31] = 0;	doodle_left_transparency_texture[36][32] = 0;	doodle_left_transparency_texture[36][33] = 0;	doodle_left_transparency_texture[36][34] = 0;	doodle_left_transparency_texture[36][35] = 0;	doodle_left_transparency_texture[36][36] = 0;	doodle_left_transparency_texture[36][37] = 0;	doodle_left_transparency_texture[36][38] = 0;	doodle_left_transparency_texture[36][39] = 0;	doodle_left_transparency_texture[36][40] = 0;	doodle_left_transparency_texture[36][41] = 0;	doodle_left_transparency_texture[36][42] = 0;	doodle_left_transparency_texture[36][43] = 0;	doodle_left_transparency_texture[36][44] = 0;	doodle_left_transparency_texture[36][45] = 0;	doodle_left_transparency_texture[36][46] = 0;	doodle_left_transparency_texture[36][47] = 0;	doodle_left_transparency_texture[36][48] = 0;	doodle_left_transparency_texture[36][49] = 0;	doodle_left_transparency_texture[36][50] = 0;	doodle_left_transparency_texture[36][51] = 0;	doodle_left_transparency_texture[36][52] = 0;	doodle_left_transparency_texture[36][53] = 0;	doodle_left_transparency_texture[36][54] = 0;	doodle_left_transparency_texture[36][55] = 0;	doodle_left_transparency_texture[36][56] = 0;	doodle_left_transparency_texture[36][57] = 0;	doodle_left_transparency_texture[36][58] = 0;	doodle_left_transparency_texture[36][59] = 0;	doodle_left_transparency_texture[36][60] = 0;	doodle_left_transparency_texture[36][61] = 0;	doodle_left_transparency_texture[36][62] = 0;	doodle_left_transparency_texture[36][63] = 0;	doodle_left_transparency_texture[36][64] = 0;	doodle_left_transparency_texture[36][65] = 0;	doodle_left_transparency_texture[36][66] = 0;	doodle_left_transparency_texture[36][67] = 0;	doodle_left_transparency_texture[36][68] = 0;	doodle_left_transparency_texture[36][69] = 0;	doodle_left_transparency_texture[36][70] = 0;	doodle_left_transparency_texture[36][71] = 0;	doodle_left_transparency_texture[36][72] = 0;	doodle_left_transparency_texture[36][73] = 0;	doodle_left_transparency_texture[36][74] = 0;	doodle_left_transparency_texture[36][75] = 0;	doodle_left_transparency_texture[36][76] = 1;	doodle_left_transparency_texture[36][77] = 1;	doodle_left_transparency_texture[36][78] = 1;	doodle_left_transparency_texture[36][79] = 1;	doodle_left_transparency_texture[37][0] = 1;	doodle_left_transparency_texture[37][1] = 1;	doodle_left_transparency_texture[37][2] = 1;	doodle_left_transparency_texture[37][3] = 1;	doodle_left_transparency_texture[37][4] = 1;	doodle_left_transparency_texture[37][5] = 1;	doodle_left_transparency_texture[37][6] = 1;	doodle_left_transparency_texture[37][7] = 1;	doodle_left_transparency_texture[37][8] = 1;	doodle_left_transparency_texture[37][9] = 1;	doodle_left_transparency_texture[37][10] = 1;	doodle_left_transparency_texture[37][11] = 1;	doodle_left_transparency_texture[37][12] = 1;	doodle_left_transparency_texture[37][13] = 1;	doodle_left_transparency_texture[37][14] = 1;	doodle_left_transparency_texture[37][15] = 1;	doodle_left_transparency_texture[37][16] = 1;	doodle_left_transparency_texture[37][17] = 1;	doodle_left_transparency_texture[37][18] = 1;	doodle_left_transparency_texture[37][19] = 1;	doodle_left_transparency_texture[37][20] = 1;	doodle_left_transparency_texture[37][21] = 1;	doodle_left_transparency_texture[37][22] = 1;	doodle_left_transparency_texture[37][23] = 1;	doodle_left_transparency_texture[37][24] = 1;	doodle_left_transparency_texture[37][25] = 1;	doodle_left_transparency_texture[37][26] = 1;	doodle_left_transparency_texture[37][27] = 1;	doodle_left_transparency_texture[37][28] = 0;	doodle_left_transparency_texture[37][29] = 0;	doodle_left_transparency_texture[37][30] = 0;	doodle_left_transparency_texture[37][31] = 0;	doodle_left_transparency_texture[37][32] = 0;	doodle_left_transparency_texture[37][33] = 0;	doodle_left_transparency_texture[37][34] = 0;	doodle_left_transparency_texture[37][35] = 0;	doodle_left_transparency_texture[37][36] = 0;	doodle_left_transparency_texture[37][37] = 0;	doodle_left_transparency_texture[37][38] = 0;	doodle_left_transparency_texture[37][39] = 0;	doodle_left_transparency_texture[37][40] = 0;	doodle_left_transparency_texture[37][41] = 0;	doodle_left_transparency_texture[37][42] = 0;	doodle_left_transparency_texture[37][43] = 0;	doodle_left_transparency_texture[37][44] = 0;	doodle_left_transparency_texture[37][45] = 0;	doodle_left_transparency_texture[37][46] = 0;	doodle_left_transparency_texture[37][47] = 0;	doodle_left_transparency_texture[37][48] = 0;	doodle_left_transparency_texture[37][49] = 0;	doodle_left_transparency_texture[37][50] = 0;	doodle_left_transparency_texture[37][51] = 0;	doodle_left_transparency_texture[37][52] = 0;	doodle_left_transparency_texture[37][53] = 0;	doodle_left_transparency_texture[37][54] = 0;	doodle_left_transparency_texture[37][55] = 0;	doodle_left_transparency_texture[37][56] = 0;	doodle_left_transparency_texture[37][57] = 0;	doodle_left_transparency_texture[37][58] = 0;	doodle_left_transparency_texture[37][59] = 0;	doodle_left_transparency_texture[37][60] = 0;	doodle_left_transparency_texture[37][61] = 0;	doodle_left_transparency_texture[37][62] = 0;	doodle_left_transparency_texture[37][63] = 0;	doodle_left_transparency_texture[37][64] = 0;	doodle_left_transparency_texture[37][65] = 0;	doodle_left_transparency_texture[37][66] = 0;	doodle_left_transparency_texture[37][67] = 0;	doodle_left_transparency_texture[37][68] = 0;	doodle_left_transparency_texture[37][69] = 0;	doodle_left_transparency_texture[37][70] = 0;	doodle_left_transparency_texture[37][71] = 0;	doodle_left_transparency_texture[37][72] = 0;	doodle_left_transparency_texture[37][73] = 0;	doodle_left_transparency_texture[37][74] = 0;	doodle_left_transparency_texture[37][75] = 0;	doodle_left_transparency_texture[37][76] = 1;	doodle_left_transparency_texture[37][77] = 1;	doodle_left_transparency_texture[37][78] = 1;	doodle_left_transparency_texture[37][79] = 1;	doodle_left_transparency_texture[38][0] = 1;	doodle_left_transparency_texture[38][1] = 1;	doodle_left_transparency_texture[38][2] = 1;	doodle_left_transparency_texture[38][3] = 1;	doodle_left_transparency_texture[38][4] = 1;	doodle_left_transparency_texture[38][5] = 1;	doodle_left_transparency_texture[38][6] = 1;	doodle_left_transparency_texture[38][7] = 1;	doodle_left_transparency_texture[38][8] = 1;	doodle_left_transparency_texture[38][9] = 1;	doodle_left_transparency_texture[38][10] = 1;	doodle_left_transparency_texture[38][11] = 1;	doodle_left_transparency_texture[38][12] = 1;	doodle_left_transparency_texture[38][13] = 1;	doodle_left_transparency_texture[38][14] = 1;	doodle_left_transparency_texture[38][15] = 1;	doodle_left_transparency_texture[38][16] = 1;	doodle_left_transparency_texture[38][17] = 1;	doodle_left_transparency_texture[38][18] = 1;	doodle_left_transparency_texture[38][19] = 1;	doodle_left_transparency_texture[38][20] = 1;	doodle_left_transparency_texture[38][21] = 1;	doodle_left_transparency_texture[38][22] = 1;	doodle_left_transparency_texture[38][23] = 1;	doodle_left_transparency_texture[38][24] = 1;	doodle_left_transparency_texture[38][25] = 1;	doodle_left_transparency_texture[38][26] = 1;	doodle_left_transparency_texture[38][27] = 1;	doodle_left_transparency_texture[38][28] = 0;	doodle_left_transparency_texture[38][29] = 0;	doodle_left_transparency_texture[38][30] = 0;	doodle_left_transparency_texture[38][31] = 0;	doodle_left_transparency_texture[38][32] = 0;	doodle_left_transparency_texture[38][33] = 0;	doodle_left_transparency_texture[38][34] = 0;	doodle_left_transparency_texture[38][35] = 0;	doodle_left_transparency_texture[38][36] = 0;	doodle_left_transparency_texture[38][37] = 0;	doodle_left_transparency_texture[38][38] = 0;	doodle_left_transparency_texture[38][39] = 0;	doodle_left_transparency_texture[38][40] = 0;	doodle_left_transparency_texture[38][41] = 0;	doodle_left_transparency_texture[38][42] = 0;	doodle_left_transparency_texture[38][43] = 0;	doodle_left_transparency_texture[38][44] = 0;	doodle_left_transparency_texture[38][45] = 0;	doodle_left_transparency_texture[38][46] = 0;	doodle_left_transparency_texture[38][47] = 0;	doodle_left_transparency_texture[38][48] = 0;	doodle_left_transparency_texture[38][49] = 0;	doodle_left_transparency_texture[38][50] = 0;	doodle_left_transparency_texture[38][51] = 0;	doodle_left_transparency_texture[38][52] = 0;	doodle_left_transparency_texture[38][53] = 0;	doodle_left_transparency_texture[38][54] = 0;	doodle_left_transparency_texture[38][55] = 0;	doodle_left_transparency_texture[38][56] = 0;	doodle_left_transparency_texture[38][57] = 0;	doodle_left_transparency_texture[38][58] = 0;	doodle_left_transparency_texture[38][59] = 0;	doodle_left_transparency_texture[38][60] = 0;	doodle_left_transparency_texture[38][61] = 0;	doodle_left_transparency_texture[38][62] = 0;	doodle_left_transparency_texture[38][63] = 0;	doodle_left_transparency_texture[38][64] = 0;	doodle_left_transparency_texture[38][65] = 0;	doodle_left_transparency_texture[38][66] = 0;	doodle_left_transparency_texture[38][67] = 0;	doodle_left_transparency_texture[38][68] = 0;	doodle_left_transparency_texture[38][69] = 0;	doodle_left_transparency_texture[38][70] = 0;	doodle_left_transparency_texture[38][71] = 0;	doodle_left_transparency_texture[38][72] = 0;	doodle_left_transparency_texture[38][73] = 0;	doodle_left_transparency_texture[38][74] = 0;	doodle_left_transparency_texture[38][75] = 0;	doodle_left_transparency_texture[38][76] = 1;	doodle_left_transparency_texture[38][77] = 1;	doodle_left_transparency_texture[38][78] = 1;	doodle_left_transparency_texture[38][79] = 1;	doodle_left_transparency_texture[39][0] = 1;	doodle_left_transparency_texture[39][1] = 1;	doodle_left_transparency_texture[39][2] = 1;	doodle_left_transparency_texture[39][3] = 1;	doodle_left_transparency_texture[39][4] = 1;	doodle_left_transparency_texture[39][5] = 1;	doodle_left_transparency_texture[39][6] = 1;	doodle_left_transparency_texture[39][7] = 1;	doodle_left_transparency_texture[39][8] = 1;	doodle_left_transparency_texture[39][9] = 1;	doodle_left_transparency_texture[39][10] = 1;	doodle_left_transparency_texture[39][11] = 1;	doodle_left_transparency_texture[39][12] = 1;	doodle_left_transparency_texture[39][13] = 1;	doodle_left_transparency_texture[39][14] = 1;	doodle_left_transparency_texture[39][15] = 1;	doodle_left_transparency_texture[39][16] = 1;	doodle_left_transparency_texture[39][17] = 1;	doodle_left_transparency_texture[39][18] = 1;	doodle_left_transparency_texture[39][19] = 1;	doodle_left_transparency_texture[39][20] = 1;	doodle_left_transparency_texture[39][21] = 1;	doodle_left_transparency_texture[39][22] = 1;	doodle_left_transparency_texture[39][23] = 1;	doodle_left_transparency_texture[39][24] = 1;	doodle_left_transparency_texture[39][25] = 1;	doodle_left_transparency_texture[39][26] = 1;	doodle_left_transparency_texture[39][27] = 1;	doodle_left_transparency_texture[39][28] = 0;	doodle_left_transparency_texture[39][29] = 0;	doodle_left_transparency_texture[39][30] = 0;	doodle_left_transparency_texture[39][31] = 0;	doodle_left_transparency_texture[39][32] = 0;	doodle_left_transparency_texture[39][33] = 0;	doodle_left_transparency_texture[39][34] = 0;	doodle_left_transparency_texture[39][35] = 0;	doodle_left_transparency_texture[39][36] = 0;	doodle_left_transparency_texture[39][37] = 0;	doodle_left_transparency_texture[39][38] = 0;	doodle_left_transparency_texture[39][39] = 0;	doodle_left_transparency_texture[39][40] = 0;	doodle_left_transparency_texture[39][41] = 0;	doodle_left_transparency_texture[39][42] = 0;	doodle_left_transparency_texture[39][43] = 0;	doodle_left_transparency_texture[39][44] = 0;	doodle_left_transparency_texture[39][45] = 0;	doodle_left_transparency_texture[39][46] = 0;	doodle_left_transparency_texture[39][47] = 0;	doodle_left_transparency_texture[39][48] = 0;	doodle_left_transparency_texture[39][49] = 0;	doodle_left_transparency_texture[39][50] = 0;	doodle_left_transparency_texture[39][51] = 0;	doodle_left_transparency_texture[39][52] = 0;	doodle_left_transparency_texture[39][53] = 0;	doodle_left_transparency_texture[39][54] = 0;	doodle_left_transparency_texture[39][55] = 0;	doodle_left_transparency_texture[39][56] = 0;	doodle_left_transparency_texture[39][57] = 0;	doodle_left_transparency_texture[39][58] = 0;	doodle_left_transparency_texture[39][59] = 0;	doodle_left_transparency_texture[39][60] = 0;	doodle_left_transparency_texture[39][61] = 0;	doodle_left_transparency_texture[39][62] = 0;	doodle_left_transparency_texture[39][63] = 0;	doodle_left_transparency_texture[39][64] = 0;	doodle_left_transparency_texture[39][65] = 0;	doodle_left_transparency_texture[39][66] = 0;	doodle_left_transparency_texture[39][67] = 0;	doodle_left_transparency_texture[39][68] = 0;	doodle_left_transparency_texture[39][69] = 0;	doodle_left_transparency_texture[39][70] = 0;	doodle_left_transparency_texture[39][71] = 0;	doodle_left_transparency_texture[39][72] = 0;	doodle_left_transparency_texture[39][73] = 0;	doodle_left_transparency_texture[39][74] = 0;	doodle_left_transparency_texture[39][75] = 0;	doodle_left_transparency_texture[39][76] = 1;	doodle_left_transparency_texture[39][77] = 1;	doodle_left_transparency_texture[39][78] = 1;	doodle_left_transparency_texture[39][79] = 1;	doodle_left_transparency_texture[40][0] = 1;	doodle_left_transparency_texture[40][1] = 1;	doodle_left_transparency_texture[40][2] = 1;	doodle_left_transparency_texture[40][3] = 1;	doodle_left_transparency_texture[40][4] = 1;	doodle_left_transparency_texture[40][5] = 1;	doodle_left_transparency_texture[40][6] = 1;	doodle_left_transparency_texture[40][7] = 1;	doodle_left_transparency_texture[40][8] = 1;	doodle_left_transparency_texture[40][9] = 1;	doodle_left_transparency_texture[40][10] = 1;	doodle_left_transparency_texture[40][11] = 1;	doodle_left_transparency_texture[40][12] = 1;	doodle_left_transparency_texture[40][13] = 1;	doodle_left_transparency_texture[40][14] = 1;	doodle_left_transparency_texture[40][15] = 1;	doodle_left_transparency_texture[40][16] = 1;	doodle_left_transparency_texture[40][17] = 1;	doodle_left_transparency_texture[40][18] = 1;	doodle_left_transparency_texture[40][19] = 1;	doodle_left_transparency_texture[40][20] = 1;	doodle_left_transparency_texture[40][21] = 1;	doodle_left_transparency_texture[40][22] = 1;	doodle_left_transparency_texture[40][23] = 1;	doodle_left_transparency_texture[40][24] = 1;	doodle_left_transparency_texture[40][25] = 1;	doodle_left_transparency_texture[40][26] = 1;	doodle_left_transparency_texture[40][27] = 1;	doodle_left_transparency_texture[40][28] = 0;	doodle_left_transparency_texture[40][29] = 0;	doodle_left_transparency_texture[40][30] = 0;	doodle_left_transparency_texture[40][31] = 0;	doodle_left_transparency_texture[40][32] = 0;	doodle_left_transparency_texture[40][33] = 0;	doodle_left_transparency_texture[40][34] = 0;	doodle_left_transparency_texture[40][35] = 0;	doodle_left_transparency_texture[40][36] = 0;	doodle_left_transparency_texture[40][37] = 0;	doodle_left_transparency_texture[40][38] = 0;	doodle_left_transparency_texture[40][39] = 0;	doodle_left_transparency_texture[40][40] = 0;	doodle_left_transparency_texture[40][41] = 0;	doodle_left_transparency_texture[40][42] = 0;	doodle_left_transparency_texture[40][43] = 0;	doodle_left_transparency_texture[40][44] = 0;	doodle_left_transparency_texture[40][45] = 0;	doodle_left_transparency_texture[40][46] = 0;	doodle_left_transparency_texture[40][47] = 0;	doodle_left_transparency_texture[40][48] = 0;	doodle_left_transparency_texture[40][49] = 0;	doodle_left_transparency_texture[40][50] = 0;	doodle_left_transparency_texture[40][51] = 0;	doodle_left_transparency_texture[40][52] = 0;	doodle_left_transparency_texture[40][53] = 0;	doodle_left_transparency_texture[40][54] = 0;	doodle_left_transparency_texture[40][55] = 0;	doodle_left_transparency_texture[40][56] = 0;	doodle_left_transparency_texture[40][57] = 0;	doodle_left_transparency_texture[40][58] = 0;	doodle_left_transparency_texture[40][59] = 0;	doodle_left_transparency_texture[40][60] = 0;	doodle_left_transparency_texture[40][61] = 0;	doodle_left_transparency_texture[40][62] = 0;	doodle_left_transparency_texture[40][63] = 0;	doodle_left_transparency_texture[40][64] = 0;	doodle_left_transparency_texture[40][65] = 0;	doodle_left_transparency_texture[40][66] = 0;	doodle_left_transparency_texture[40][67] = 0;	doodle_left_transparency_texture[40][68] = 0;	doodle_left_transparency_texture[40][69] = 0;	doodle_left_transparency_texture[40][70] = 0;	doodle_left_transparency_texture[40][71] = 0;	doodle_left_transparency_texture[40][72] = 0;	doodle_left_transparency_texture[40][73] = 0;	doodle_left_transparency_texture[40][74] = 0;	doodle_left_transparency_texture[40][75] = 0;	doodle_left_transparency_texture[40][76] = 1;	doodle_left_transparency_texture[40][77] = 1;	doodle_left_transparency_texture[40][78] = 1;	doodle_left_transparency_texture[40][79] = 1;	doodle_left_transparency_texture[41][0] = 1;	doodle_left_transparency_texture[41][1] = 1;	doodle_left_transparency_texture[41][2] = 1;	doodle_left_transparency_texture[41][3] = 1;	doodle_left_transparency_texture[41][4] = 1;	doodle_left_transparency_texture[41][5] = 1;	doodle_left_transparency_texture[41][6] = 1;	doodle_left_transparency_texture[41][7] = 1;	doodle_left_transparency_texture[41][8] = 1;	doodle_left_transparency_texture[41][9] = 1;	doodle_left_transparency_texture[41][10] = 1;	doodle_left_transparency_texture[41][11] = 1;	doodle_left_transparency_texture[41][12] = 1;	doodle_left_transparency_texture[41][13] = 1;	doodle_left_transparency_texture[41][14] = 1;	doodle_left_transparency_texture[41][15] = 1;	doodle_left_transparency_texture[41][16] = 1;	doodle_left_transparency_texture[41][17] = 1;	doodle_left_transparency_texture[41][18] = 1;	doodle_left_transparency_texture[41][19] = 1;	doodle_left_transparency_texture[41][20] = 1;	doodle_left_transparency_texture[41][21] = 1;	doodle_left_transparency_texture[41][22] = 1;	doodle_left_transparency_texture[41][23] = 1;	doodle_left_transparency_texture[41][24] = 1;	doodle_left_transparency_texture[41][25] = 1;	doodle_left_transparency_texture[41][26] = 1;	doodle_left_transparency_texture[41][27] = 1;	doodle_left_transparency_texture[41][28] = 0;	doodle_left_transparency_texture[41][29] = 0;	doodle_left_transparency_texture[41][30] = 0;	doodle_left_transparency_texture[41][31] = 0;	doodle_left_transparency_texture[41][32] = 0;	doodle_left_transparency_texture[41][33] = 0;	doodle_left_transparency_texture[41][34] = 0;	doodle_left_transparency_texture[41][35] = 0;	doodle_left_transparency_texture[41][36] = 0;	doodle_left_transparency_texture[41][37] = 0;	doodle_left_transparency_texture[41][38] = 0;	doodle_left_transparency_texture[41][39] = 0;	doodle_left_transparency_texture[41][40] = 0;	doodle_left_transparency_texture[41][41] = 0;	doodle_left_transparency_texture[41][42] = 0;	doodle_left_transparency_texture[41][43] = 0;	doodle_left_transparency_texture[41][44] = 0;	doodle_left_transparency_texture[41][45] = 0;	doodle_left_transparency_texture[41][46] = 0;	doodle_left_transparency_texture[41][47] = 0;	doodle_left_transparency_texture[41][48] = 0;	doodle_left_transparency_texture[41][49] = 0;	doodle_left_transparency_texture[41][50] = 0;	doodle_left_transparency_texture[41][51] = 0;	doodle_left_transparency_texture[41][52] = 0;	doodle_left_transparency_texture[41][53] = 0;	doodle_left_transparency_texture[41][54] = 0;	doodle_left_transparency_texture[41][55] = 0;	doodle_left_transparency_texture[41][56] = 0;	doodle_left_transparency_texture[41][57] = 0;	doodle_left_transparency_texture[41][58] = 0;	doodle_left_transparency_texture[41][59] = 0;	doodle_left_transparency_texture[41][60] = 0;	doodle_left_transparency_texture[41][61] = 0;	doodle_left_transparency_texture[41][62] = 0;	doodle_left_transparency_texture[41][63] = 0;	doodle_left_transparency_texture[41][64] = 0;	doodle_left_transparency_texture[41][65] = 0;	doodle_left_transparency_texture[41][66] = 0;	doodle_left_transparency_texture[41][67] = 0;	doodle_left_transparency_texture[41][68] = 0;	doodle_left_transparency_texture[41][69] = 0;	doodle_left_transparency_texture[41][70] = 0;	doodle_left_transparency_texture[41][71] = 0;	doodle_left_transparency_texture[41][72] = 0;	doodle_left_transparency_texture[41][73] = 0;	doodle_left_transparency_texture[41][74] = 0;	doodle_left_transparency_texture[41][75] = 0;	doodle_left_transparency_texture[41][76] = 1;	doodle_left_transparency_texture[41][77] = 1;	doodle_left_transparency_texture[41][78] = 1;	doodle_left_transparency_texture[41][79] = 1;	doodle_left_transparency_texture[42][0] = 1;	doodle_left_transparency_texture[42][1] = 1;	doodle_left_transparency_texture[42][2] = 1;	doodle_left_transparency_texture[42][3] = 1;	doodle_left_transparency_texture[42][4] = 1;	doodle_left_transparency_texture[42][5] = 1;	doodle_left_transparency_texture[42][6] = 1;	doodle_left_transparency_texture[42][7] = 1;	doodle_left_transparency_texture[42][8] = 1;	doodle_left_transparency_texture[42][9] = 1;	doodle_left_transparency_texture[42][10] = 1;	doodle_left_transparency_texture[42][11] = 1;	doodle_left_transparency_texture[42][12] = 1;	doodle_left_transparency_texture[42][13] = 1;	doodle_left_transparency_texture[42][14] = 1;	doodle_left_transparency_texture[42][15] = 1;	doodle_left_transparency_texture[42][16] = 1;	doodle_left_transparency_texture[42][17] = 1;	doodle_left_transparency_texture[42][18] = 1;	doodle_left_transparency_texture[42][19] = 1;	doodle_left_transparency_texture[42][20] = 1;	doodle_left_transparency_texture[42][21] = 1;	doodle_left_transparency_texture[42][22] = 1;	doodle_left_transparency_texture[42][23] = 1;	doodle_left_transparency_texture[42][24] = 1;	doodle_left_transparency_texture[42][25] = 1;	doodle_left_transparency_texture[42][26] = 1;	doodle_left_transparency_texture[42][27] = 1;	doodle_left_transparency_texture[42][28] = 0;	doodle_left_transparency_texture[42][29] = 0;	doodle_left_transparency_texture[42][30] = 0;	doodle_left_transparency_texture[42][31] = 0;	doodle_left_transparency_texture[42][32] = 0;	doodle_left_transparency_texture[42][33] = 0;	doodle_left_transparency_texture[42][34] = 0;	doodle_left_transparency_texture[42][35] = 0;	doodle_left_transparency_texture[42][36] = 0;	doodle_left_transparency_texture[42][37] = 0;	doodle_left_transparency_texture[42][38] = 0;	doodle_left_transparency_texture[42][39] = 0;	doodle_left_transparency_texture[42][40] = 0;	doodle_left_transparency_texture[42][41] = 0;	doodle_left_transparency_texture[42][42] = 0;	doodle_left_transparency_texture[42][43] = 0;	doodle_left_transparency_texture[42][44] = 0;	doodle_left_transparency_texture[42][45] = 0;	doodle_left_transparency_texture[42][46] = 0;	doodle_left_transparency_texture[42][47] = 0;	doodle_left_transparency_texture[42][48] = 0;	doodle_left_transparency_texture[42][49] = 0;	doodle_left_transparency_texture[42][50] = 0;	doodle_left_transparency_texture[42][51] = 0;	doodle_left_transparency_texture[42][52] = 0;	doodle_left_transparency_texture[42][53] = 0;	doodle_left_transparency_texture[42][54] = 0;	doodle_left_transparency_texture[42][55] = 0;	doodle_left_transparency_texture[42][56] = 0;	doodle_left_transparency_texture[42][57] = 0;	doodle_left_transparency_texture[42][58] = 0;	doodle_left_transparency_texture[42][59] = 0;	doodle_left_transparency_texture[42][60] = 0;	doodle_left_transparency_texture[42][61] = 0;	doodle_left_transparency_texture[42][62] = 0;	doodle_left_transparency_texture[42][63] = 0;	doodle_left_transparency_texture[42][64] = 0;	doodle_left_transparency_texture[42][65] = 0;	doodle_left_transparency_texture[42][66] = 0;	doodle_left_transparency_texture[42][67] = 0;	doodle_left_transparency_texture[42][68] = 0;	doodle_left_transparency_texture[42][69] = 0;	doodle_left_transparency_texture[42][70] = 0;	doodle_left_transparency_texture[42][71] = 0;	doodle_left_transparency_texture[42][72] = 0;	doodle_left_transparency_texture[42][73] = 0;	doodle_left_transparency_texture[42][74] = 0;	doodle_left_transparency_texture[42][75] = 0;	doodle_left_transparency_texture[42][76] = 1;	doodle_left_transparency_texture[42][77] = 1;	doodle_left_transparency_texture[42][78] = 1;	doodle_left_transparency_texture[42][79] = 1;	doodle_left_transparency_texture[43][0] = 1;	doodle_left_transparency_texture[43][1] = 1;	doodle_left_transparency_texture[43][2] = 1;	doodle_left_transparency_texture[43][3] = 1;	doodle_left_transparency_texture[43][4] = 1;	doodle_left_transparency_texture[43][5] = 1;	doodle_left_transparency_texture[43][6] = 1;	doodle_left_transparency_texture[43][7] = 1;	doodle_left_transparency_texture[43][8] = 1;	doodle_left_transparency_texture[43][9] = 1;	doodle_left_transparency_texture[43][10] = 1;	doodle_left_transparency_texture[43][11] = 1;	doodle_left_transparency_texture[43][12] = 1;	doodle_left_transparency_texture[43][13] = 1;	doodle_left_transparency_texture[43][14] = 1;	doodle_left_transparency_texture[43][15] = 1;	doodle_left_transparency_texture[43][16] = 1;	doodle_left_transparency_texture[43][17] = 1;	doodle_left_transparency_texture[43][18] = 1;	doodle_left_transparency_texture[43][19] = 1;	doodle_left_transparency_texture[43][20] = 1;	doodle_left_transparency_texture[43][21] = 1;	doodle_left_transparency_texture[43][22] = 1;	doodle_left_transparency_texture[43][23] = 1;	doodle_left_transparency_texture[43][24] = 1;	doodle_left_transparency_texture[43][25] = 1;	doodle_left_transparency_texture[43][26] = 1;	doodle_left_transparency_texture[43][27] = 1;	doodle_left_transparency_texture[43][28] = 0;	doodle_left_transparency_texture[43][29] = 0;	doodle_left_transparency_texture[43][30] = 0;	doodle_left_transparency_texture[43][31] = 0;	doodle_left_transparency_texture[43][32] = 0;	doodle_left_transparency_texture[43][33] = 0;	doodle_left_transparency_texture[43][34] = 0;	doodle_left_transparency_texture[43][35] = 0;	doodle_left_transparency_texture[43][36] = 0;	doodle_left_transparency_texture[43][37] = 0;	doodle_left_transparency_texture[43][38] = 0;	doodle_left_transparency_texture[43][39] = 0;	doodle_left_transparency_texture[43][40] = 0;	doodle_left_transparency_texture[43][41] = 0;	doodle_left_transparency_texture[43][42] = 0;	doodle_left_transparency_texture[43][43] = 0;	doodle_left_transparency_texture[43][44] = 0;	doodle_left_transparency_texture[43][45] = 0;	doodle_left_transparency_texture[43][46] = 0;	doodle_left_transparency_texture[43][47] = 0;	doodle_left_transparency_texture[43][48] = 0;	doodle_left_transparency_texture[43][49] = 0;	doodle_left_transparency_texture[43][50] = 0;	doodle_left_transparency_texture[43][51] = 0;	doodle_left_transparency_texture[43][52] = 0;	doodle_left_transparency_texture[43][53] = 0;	doodle_left_transparency_texture[43][54] = 0;	doodle_left_transparency_texture[43][55] = 0;	doodle_left_transparency_texture[43][56] = 0;	doodle_left_transparency_texture[43][57] = 0;	doodle_left_transparency_texture[43][58] = 0;	doodle_left_transparency_texture[43][59] = 0;	doodle_left_transparency_texture[43][60] = 0;	doodle_left_transparency_texture[43][61] = 0;	doodle_left_transparency_texture[43][62] = 0;	doodle_left_transparency_texture[43][63] = 0;	doodle_left_transparency_texture[43][64] = 0;	doodle_left_transparency_texture[43][65] = 0;	doodle_left_transparency_texture[43][66] = 0;	doodle_left_transparency_texture[43][67] = 0;	doodle_left_transparency_texture[43][68] = 0;	doodle_left_transparency_texture[43][69] = 0;	doodle_left_transparency_texture[43][70] = 0;	doodle_left_transparency_texture[43][71] = 0;	doodle_left_transparency_texture[43][72] = 0;	doodle_left_transparency_texture[43][73] = 0;	doodle_left_transparency_texture[43][74] = 0;	doodle_left_transparency_texture[43][75] = 0;	doodle_left_transparency_texture[43][76] = 1;	doodle_left_transparency_texture[43][77] = 1;	doodle_left_transparency_texture[43][78] = 1;	doodle_left_transparency_texture[43][79] = 1;	doodle_left_transparency_texture[44][0] = 1;	doodle_left_transparency_texture[44][1] = 1;	doodle_left_transparency_texture[44][2] = 1;	doodle_left_transparency_texture[44][3] = 1;	doodle_left_transparency_texture[44][4] = 1;	doodle_left_transparency_texture[44][5] = 1;	doodle_left_transparency_texture[44][6] = 1;	doodle_left_transparency_texture[44][7] = 1;	doodle_left_transparency_texture[44][8] = 1;	doodle_left_transparency_texture[44][9] = 1;	doodle_left_transparency_texture[44][10] = 1;	doodle_left_transparency_texture[44][11] = 1;	doodle_left_transparency_texture[44][12] = 1;	doodle_left_transparency_texture[44][13] = 1;	doodle_left_transparency_texture[44][14] = 1;	doodle_left_transparency_texture[44][15] = 1;	doodle_left_transparency_texture[44][16] = 1;	doodle_left_transparency_texture[44][17] = 1;	doodle_left_transparency_texture[44][18] = 1;	doodle_left_transparency_texture[44][19] = 1;	doodle_left_transparency_texture[44][20] = 1;	doodle_left_transparency_texture[44][21] = 1;	doodle_left_transparency_texture[44][22] = 1;	doodle_left_transparency_texture[44][23] = 1;	doodle_left_transparency_texture[44][24] = 1;	doodle_left_transparency_texture[44][25] = 1;	doodle_left_transparency_texture[44][26] = 1;	doodle_left_transparency_texture[44][27] = 1;	doodle_left_transparency_texture[44][28] = 0;	doodle_left_transparency_texture[44][29] = 0;	doodle_left_transparency_texture[44][30] = 0;	doodle_left_transparency_texture[44][31] = 0;	doodle_left_transparency_texture[44][32] = 0;	doodle_left_transparency_texture[44][33] = 0;	doodle_left_transparency_texture[44][34] = 0;	doodle_left_transparency_texture[44][35] = 0;	doodle_left_transparency_texture[44][36] = 0;	doodle_left_transparency_texture[44][37] = 0;	doodle_left_transparency_texture[44][38] = 0;	doodle_left_transparency_texture[44][39] = 0;	doodle_left_transparency_texture[44][40] = 0;	doodle_left_transparency_texture[44][41] = 0;	doodle_left_transparency_texture[44][42] = 0;	doodle_left_transparency_texture[44][43] = 0;	doodle_left_transparency_texture[44][44] = 0;	doodle_left_transparency_texture[44][45] = 0;	doodle_left_transparency_texture[44][46] = 0;	doodle_left_transparency_texture[44][47] = 0;	doodle_left_transparency_texture[44][48] = 0;	doodle_left_transparency_texture[44][49] = 0;	doodle_left_transparency_texture[44][50] = 0;	doodle_left_transparency_texture[44][51] = 0;	doodle_left_transparency_texture[44][52] = 0;	doodle_left_transparency_texture[44][53] = 0;	doodle_left_transparency_texture[44][54] = 0;	doodle_left_transparency_texture[44][55] = 0;	doodle_left_transparency_texture[44][56] = 0;	doodle_left_transparency_texture[44][57] = 0;	doodle_left_transparency_texture[44][58] = 0;	doodle_left_transparency_texture[44][59] = 0;	doodle_left_transparency_texture[44][60] = 0;	doodle_left_transparency_texture[44][61] = 0;	doodle_left_transparency_texture[44][62] = 0;	doodle_left_transparency_texture[44][63] = 0;	doodle_left_transparency_texture[44][64] = 0;	doodle_left_transparency_texture[44][65] = 0;	doodle_left_transparency_texture[44][66] = 0;	doodle_left_transparency_texture[44][67] = 0;	doodle_left_transparency_texture[44][68] = 0;	doodle_left_transparency_texture[44][69] = 0;	doodle_left_transparency_texture[44][70] = 0;	doodle_left_transparency_texture[44][71] = 0;	doodle_left_transparency_texture[44][72] = 0;	doodle_left_transparency_texture[44][73] = 0;	doodle_left_transparency_texture[44][74] = 0;	doodle_left_transparency_texture[44][75] = 0;	doodle_left_transparency_texture[44][76] = 1;	doodle_left_transparency_texture[44][77] = 1;	doodle_left_transparency_texture[44][78] = 1;	doodle_left_transparency_texture[44][79] = 1;	doodle_left_transparency_texture[45][0] = 1;	doodle_left_transparency_texture[45][1] = 1;	doodle_left_transparency_texture[45][2] = 1;	doodle_left_transparency_texture[45][3] = 1;	doodle_left_transparency_texture[45][4] = 1;	doodle_left_transparency_texture[45][5] = 1;	doodle_left_transparency_texture[45][6] = 1;	doodle_left_transparency_texture[45][7] = 1;	doodle_left_transparency_texture[45][8] = 1;	doodle_left_transparency_texture[45][9] = 1;	doodle_left_transparency_texture[45][10] = 1;	doodle_left_transparency_texture[45][11] = 1;	doodle_left_transparency_texture[45][12] = 1;	doodle_left_transparency_texture[45][13] = 1;	doodle_left_transparency_texture[45][14] = 1;	doodle_left_transparency_texture[45][15] = 1;	doodle_left_transparency_texture[45][16] = 1;	doodle_left_transparency_texture[45][17] = 1;	doodle_left_transparency_texture[45][18] = 1;	doodle_left_transparency_texture[45][19] = 1;	doodle_left_transparency_texture[45][20] = 1;	doodle_left_transparency_texture[45][21] = 1;	doodle_left_transparency_texture[45][22] = 1;	doodle_left_transparency_texture[45][23] = 1;	doodle_left_transparency_texture[45][24] = 1;	doodle_left_transparency_texture[45][25] = 1;	doodle_left_transparency_texture[45][26] = 1;	doodle_left_transparency_texture[45][27] = 1;	doodle_left_transparency_texture[45][28] = 0;	doodle_left_transparency_texture[45][29] = 0;	doodle_left_transparency_texture[45][30] = 0;	doodle_left_transparency_texture[45][31] = 0;	doodle_left_transparency_texture[45][32] = 0;	doodle_left_transparency_texture[45][33] = 0;	doodle_left_transparency_texture[45][34] = 0;	doodle_left_transparency_texture[45][35] = 0;	doodle_left_transparency_texture[45][36] = 0;	doodle_left_transparency_texture[45][37] = 0;	doodle_left_transparency_texture[45][38] = 0;	doodle_left_transparency_texture[45][39] = 0;	doodle_left_transparency_texture[45][40] = 0;	doodle_left_transparency_texture[45][41] = 0;	doodle_left_transparency_texture[45][42] = 0;	doodle_left_transparency_texture[45][43] = 0;	doodle_left_transparency_texture[45][44] = 0;	doodle_left_transparency_texture[45][45] = 0;	doodle_left_transparency_texture[45][46] = 0;	doodle_left_transparency_texture[45][47] = 0;	doodle_left_transparency_texture[45][48] = 0;	doodle_left_transparency_texture[45][49] = 0;	doodle_left_transparency_texture[45][50] = 0;	doodle_left_transparency_texture[45][51] = 0;	doodle_left_transparency_texture[45][52] = 0;	doodle_left_transparency_texture[45][53] = 0;	doodle_left_transparency_texture[45][54] = 0;	doodle_left_transparency_texture[45][55] = 0;	doodle_left_transparency_texture[45][56] = 0;	doodle_left_transparency_texture[45][57] = 0;	doodle_left_transparency_texture[45][58] = 0;	doodle_left_transparency_texture[45][59] = 0;	doodle_left_transparency_texture[45][60] = 0;	doodle_left_transparency_texture[45][61] = 0;	doodle_left_transparency_texture[45][62] = 0;	doodle_left_transparency_texture[45][63] = 0;	doodle_left_transparency_texture[45][64] = 0;	doodle_left_transparency_texture[45][65] = 0;	doodle_left_transparency_texture[45][66] = 0;	doodle_left_transparency_texture[45][67] = 0;	doodle_left_transparency_texture[45][68] = 0;	doodle_left_transparency_texture[45][69] = 0;	doodle_left_transparency_texture[45][70] = 0;	doodle_left_transparency_texture[45][71] = 0;	doodle_left_transparency_texture[45][72] = 0;	doodle_left_transparency_texture[45][73] = 0;	doodle_left_transparency_texture[45][74] = 0;	doodle_left_transparency_texture[45][75] = 0;	doodle_left_transparency_texture[45][76] = 1;	doodle_left_transparency_texture[45][77] = 1;	doodle_left_transparency_texture[45][78] = 1;	doodle_left_transparency_texture[45][79] = 1;	doodle_left_transparency_texture[46][0] = 1;	doodle_left_transparency_texture[46][1] = 1;	doodle_left_transparency_texture[46][2] = 1;	doodle_left_transparency_texture[46][3] = 1;	doodle_left_transparency_texture[46][4] = 1;	doodle_left_transparency_texture[46][5] = 1;	doodle_left_transparency_texture[46][6] = 1;	doodle_left_transparency_texture[46][7] = 1;	doodle_left_transparency_texture[46][8] = 1;	doodle_left_transparency_texture[46][9] = 1;	doodle_left_transparency_texture[46][10] = 1;	doodle_left_transparency_texture[46][11] = 1;	doodle_left_transparency_texture[46][12] = 1;	doodle_left_transparency_texture[46][13] = 1;	doodle_left_transparency_texture[46][14] = 1;	doodle_left_transparency_texture[46][15] = 1;	doodle_left_transparency_texture[46][16] = 1;	doodle_left_transparency_texture[46][17] = 1;	doodle_left_transparency_texture[46][18] = 1;	doodle_left_transparency_texture[46][19] = 1;	doodle_left_transparency_texture[46][20] = 1;	doodle_left_transparency_texture[46][21] = 1;	doodle_left_transparency_texture[46][22] = 1;	doodle_left_transparency_texture[46][23] = 1;	doodle_left_transparency_texture[46][24] = 1;	doodle_left_transparency_texture[46][25] = 1;	doodle_left_transparency_texture[46][26] = 1;	doodle_left_transparency_texture[46][27] = 1;	doodle_left_transparency_texture[46][28] = 0;	doodle_left_transparency_texture[46][29] = 0;	doodle_left_transparency_texture[46][30] = 0;	doodle_left_transparency_texture[46][31] = 0;	doodle_left_transparency_texture[46][32] = 0;	doodle_left_transparency_texture[46][33] = 0;	doodle_left_transparency_texture[46][34] = 0;	doodle_left_transparency_texture[46][35] = 0;	doodle_left_transparency_texture[46][36] = 0;	doodle_left_transparency_texture[46][37] = 0;	doodle_left_transparency_texture[46][38] = 0;	doodle_left_transparency_texture[46][39] = 0;	doodle_left_transparency_texture[46][40] = 0;	doodle_left_transparency_texture[46][41] = 0;	doodle_left_transparency_texture[46][42] = 0;	doodle_left_transparency_texture[46][43] = 0;	doodle_left_transparency_texture[46][44] = 0;	doodle_left_transparency_texture[46][45] = 0;	doodle_left_transparency_texture[46][46] = 0;	doodle_left_transparency_texture[46][47] = 0;	doodle_left_transparency_texture[46][48] = 0;	doodle_left_transparency_texture[46][49] = 0;	doodle_left_transparency_texture[46][50] = 0;	doodle_left_transparency_texture[46][51] = 0;	doodle_left_transparency_texture[46][52] = 0;	doodle_left_transparency_texture[46][53] = 0;	doodle_left_transparency_texture[46][54] = 0;	doodle_left_transparency_texture[46][55] = 0;	doodle_left_transparency_texture[46][56] = 0;	doodle_left_transparency_texture[46][57] = 0;	doodle_left_transparency_texture[46][58] = 0;	doodle_left_transparency_texture[46][59] = 0;	doodle_left_transparency_texture[46][60] = 0;	doodle_left_transparency_texture[46][61] = 0;	doodle_left_transparency_texture[46][62] = 0;	doodle_left_transparency_texture[46][63] = 0;	doodle_left_transparency_texture[46][64] = 0;	doodle_left_transparency_texture[46][65] = 0;	doodle_left_transparency_texture[46][66] = 0;	doodle_left_transparency_texture[46][67] = 0;	doodle_left_transparency_texture[46][68] = 0;	doodle_left_transparency_texture[46][69] = 0;	doodle_left_transparency_texture[46][70] = 0;	doodle_left_transparency_texture[46][71] = 0;	doodle_left_transparency_texture[46][72] = 0;	doodle_left_transparency_texture[46][73] = 0;	doodle_left_transparency_texture[46][74] = 0;	doodle_left_transparency_texture[46][75] = 0;	doodle_left_transparency_texture[46][76] = 1;	doodle_left_transparency_texture[46][77] = 1;	doodle_left_transparency_texture[46][78] = 1;	doodle_left_transparency_texture[46][79] = 1;	doodle_left_transparency_texture[47][0] = 1;	doodle_left_transparency_texture[47][1] = 1;	doodle_left_transparency_texture[47][2] = 1;	doodle_left_transparency_texture[47][3] = 1;	doodle_left_transparency_texture[47][4] = 1;	doodle_left_transparency_texture[47][5] = 1;	doodle_left_transparency_texture[47][6] = 1;	doodle_left_transparency_texture[47][7] = 1;	doodle_left_transparency_texture[47][8] = 1;	doodle_left_transparency_texture[47][9] = 1;	doodle_left_transparency_texture[47][10] = 1;	doodle_left_transparency_texture[47][11] = 1;	doodle_left_transparency_texture[47][12] = 1;	doodle_left_transparency_texture[47][13] = 1;	doodle_left_transparency_texture[47][14] = 1;	doodle_left_transparency_texture[47][15] = 1;	doodle_left_transparency_texture[47][16] = 1;	doodle_left_transparency_texture[47][17] = 1;	doodle_left_transparency_texture[47][18] = 1;	doodle_left_transparency_texture[47][19] = 1;	doodle_left_transparency_texture[47][20] = 1;	doodle_left_transparency_texture[47][21] = 1;	doodle_left_transparency_texture[47][22] = 1;	doodle_left_transparency_texture[47][23] = 1;	doodle_left_transparency_texture[47][24] = 1;	doodle_left_transparency_texture[47][25] = 1;	doodle_left_transparency_texture[47][26] = 1;	doodle_left_transparency_texture[47][27] = 1;	doodle_left_transparency_texture[47][28] = 0;	doodle_left_transparency_texture[47][29] = 0;	doodle_left_transparency_texture[47][30] = 0;	doodle_left_transparency_texture[47][31] = 0;	doodle_left_transparency_texture[47][32] = 0;	doodle_left_transparency_texture[47][33] = 0;	doodle_left_transparency_texture[47][34] = 0;	doodle_left_transparency_texture[47][35] = 0;	doodle_left_transparency_texture[47][36] = 0;	doodle_left_transparency_texture[47][37] = 0;	doodle_left_transparency_texture[47][38] = 0;	doodle_left_transparency_texture[47][39] = 0;	doodle_left_transparency_texture[47][40] = 0;	doodle_left_transparency_texture[47][41] = 0;	doodle_left_transparency_texture[47][42] = 0;	doodle_left_transparency_texture[47][43] = 0;	doodle_left_transparency_texture[47][44] = 0;	doodle_left_transparency_texture[47][45] = 0;	doodle_left_transparency_texture[47][46] = 0;	doodle_left_transparency_texture[47][47] = 0;	doodle_left_transparency_texture[47][48] = 0;	doodle_left_transparency_texture[47][49] = 0;	doodle_left_transparency_texture[47][50] = 0;	doodle_left_transparency_texture[47][51] = 0;	doodle_left_transparency_texture[47][52] = 0;	doodle_left_transparency_texture[47][53] = 0;	doodle_left_transparency_texture[47][54] = 0;	doodle_left_transparency_texture[47][55] = 0;	doodle_left_transparency_texture[47][56] = 0;	doodle_left_transparency_texture[47][57] = 0;	doodle_left_transparency_texture[47][58] = 0;	doodle_left_transparency_texture[47][59] = 0;	doodle_left_transparency_texture[47][60] = 0;	doodle_left_transparency_texture[47][61] = 0;	doodle_left_transparency_texture[47][62] = 0;	doodle_left_transparency_texture[47][63] = 0;	doodle_left_transparency_texture[47][64] = 0;	doodle_left_transparency_texture[47][65] = 0;	doodle_left_transparency_texture[47][66] = 0;	doodle_left_transparency_texture[47][67] = 0;	doodle_left_transparency_texture[47][68] = 0;	doodle_left_transparency_texture[47][69] = 0;	doodle_left_transparency_texture[47][70] = 0;	doodle_left_transparency_texture[47][71] = 0;	doodle_left_transparency_texture[47][72] = 0;	doodle_left_transparency_texture[47][73] = 0;	doodle_left_transparency_texture[47][74] = 0;	doodle_left_transparency_texture[47][75] = 0;	doodle_left_transparency_texture[47][76] = 1;	doodle_left_transparency_texture[47][77] = 1;	doodle_left_transparency_texture[47][78] = 1;	doodle_left_transparency_texture[47][79] = 1;	doodle_left_transparency_texture[48][0] = 1;	doodle_left_transparency_texture[48][1] = 1;	doodle_left_transparency_texture[48][2] = 1;	doodle_left_transparency_texture[48][3] = 1;	doodle_left_transparency_texture[48][4] = 1;	doodle_left_transparency_texture[48][5] = 1;	doodle_left_transparency_texture[48][6] = 1;	doodle_left_transparency_texture[48][7] = 1;	doodle_left_transparency_texture[48][8] = 1;	doodle_left_transparency_texture[48][9] = 1;	doodle_left_transparency_texture[48][10] = 1;	doodle_left_transparency_texture[48][11] = 1;	doodle_left_transparency_texture[48][12] = 1;	doodle_left_transparency_texture[48][13] = 1;	doodle_left_transparency_texture[48][14] = 1;	doodle_left_transparency_texture[48][15] = 1;	doodle_left_transparency_texture[48][16] = 1;	doodle_left_transparency_texture[48][17] = 1;	doodle_left_transparency_texture[48][18] = 1;	doodle_left_transparency_texture[48][19] = 1;	doodle_left_transparency_texture[48][20] = 1;	doodle_left_transparency_texture[48][21] = 1;	doodle_left_transparency_texture[48][22] = 1;	doodle_left_transparency_texture[48][23] = 1;	doodle_left_transparency_texture[48][24] = 1;	doodle_left_transparency_texture[48][25] = 1;	doodle_left_transparency_texture[48][26] = 1;	doodle_left_transparency_texture[48][27] = 1;	doodle_left_transparency_texture[48][28] = 0;	doodle_left_transparency_texture[48][29] = 0;	doodle_left_transparency_texture[48][30] = 0;	doodle_left_transparency_texture[48][31] = 0;	doodle_left_transparency_texture[48][32] = 0;	doodle_left_transparency_texture[48][33] = 0;	doodle_left_transparency_texture[48][34] = 0;	doodle_left_transparency_texture[48][35] = 0;	doodle_left_transparency_texture[48][36] = 0;	doodle_left_transparency_texture[48][37] = 0;	doodle_left_transparency_texture[48][38] = 0;	doodle_left_transparency_texture[48][39] = 0;	doodle_left_transparency_texture[48][40] = 0;	doodle_left_transparency_texture[48][41] = 0;	doodle_left_transparency_texture[48][42] = 0;	doodle_left_transparency_texture[48][43] = 0;	doodle_left_transparency_texture[48][44] = 0;	doodle_left_transparency_texture[48][45] = 0;	doodle_left_transparency_texture[48][46] = 0;	doodle_left_transparency_texture[48][47] = 0;	doodle_left_transparency_texture[48][48] = 0;	doodle_left_transparency_texture[48][49] = 0;	doodle_left_transparency_texture[48][50] = 0;	doodle_left_transparency_texture[48][51] = 0;	doodle_left_transparency_texture[48][52] = 0;	doodle_left_transparency_texture[48][53] = 0;	doodle_left_transparency_texture[48][54] = 0;	doodle_left_transparency_texture[48][55] = 0;	doodle_left_transparency_texture[48][56] = 0;	doodle_left_transparency_texture[48][57] = 0;	doodle_left_transparency_texture[48][58] = 0;	doodle_left_transparency_texture[48][59] = 0;	doodle_left_transparency_texture[48][60] = 0;	doodle_left_transparency_texture[48][61] = 0;	doodle_left_transparency_texture[48][62] = 0;	doodle_left_transparency_texture[48][63] = 0;	doodle_left_transparency_texture[48][64] = 0;	doodle_left_transparency_texture[48][65] = 0;	doodle_left_transparency_texture[48][66] = 0;	doodle_left_transparency_texture[48][67] = 0;	doodle_left_transparency_texture[48][68] = 0;	doodle_left_transparency_texture[48][69] = 0;	doodle_left_transparency_texture[48][70] = 0;	doodle_left_transparency_texture[48][71] = 0;	doodle_left_transparency_texture[48][72] = 0;	doodle_left_transparency_texture[48][73] = 0;	doodle_left_transparency_texture[48][74] = 0;	doodle_left_transparency_texture[48][75] = 0;	doodle_left_transparency_texture[48][76] = 1;	doodle_left_transparency_texture[48][77] = 1;	doodle_left_transparency_texture[48][78] = 1;	doodle_left_transparency_texture[48][79] = 1;	doodle_left_transparency_texture[49][0] = 1;	doodle_left_transparency_texture[49][1] = 1;	doodle_left_transparency_texture[49][2] = 1;	doodle_left_transparency_texture[49][3] = 1;	doodle_left_transparency_texture[49][4] = 1;	doodle_left_transparency_texture[49][5] = 1;	doodle_left_transparency_texture[49][6] = 1;	doodle_left_transparency_texture[49][7] = 1;	doodle_left_transparency_texture[49][8] = 1;	doodle_left_transparency_texture[49][9] = 1;	doodle_left_transparency_texture[49][10] = 1;	doodle_left_transparency_texture[49][11] = 1;	doodle_left_transparency_texture[49][12] = 1;	doodle_left_transparency_texture[49][13] = 1;	doodle_left_transparency_texture[49][14] = 1;	doodle_left_transparency_texture[49][15] = 1;	doodle_left_transparency_texture[49][16] = 1;	doodle_left_transparency_texture[49][17] = 1;	doodle_left_transparency_texture[49][18] = 1;	doodle_left_transparency_texture[49][19] = 1;	doodle_left_transparency_texture[49][20] = 1;	doodle_left_transparency_texture[49][21] = 1;	doodle_left_transparency_texture[49][22] = 1;	doodle_left_transparency_texture[49][23] = 1;	doodle_left_transparency_texture[49][24] = 1;	doodle_left_transparency_texture[49][25] = 1;	doodle_left_transparency_texture[49][26] = 1;	doodle_left_transparency_texture[49][27] = 1;	doodle_left_transparency_texture[49][28] = 0;	doodle_left_transparency_texture[49][29] = 0;	doodle_left_transparency_texture[49][30] = 0;	doodle_left_transparency_texture[49][31] = 0;	doodle_left_transparency_texture[49][32] = 0;	doodle_left_transparency_texture[49][33] = 0;	doodle_left_transparency_texture[49][34] = 0;	doodle_left_transparency_texture[49][35] = 0;	doodle_left_transparency_texture[49][36] = 0;	doodle_left_transparency_texture[49][37] = 0;	doodle_left_transparency_texture[49][38] = 0;	doodle_left_transparency_texture[49][39] = 0;	doodle_left_transparency_texture[49][40] = 0;	doodle_left_transparency_texture[49][41] = 0;	doodle_left_transparency_texture[49][42] = 0;	doodle_left_transparency_texture[49][43] = 0;	doodle_left_transparency_texture[49][44] = 0;	doodle_left_transparency_texture[49][45] = 0;	doodle_left_transparency_texture[49][46] = 0;	doodle_left_transparency_texture[49][47] = 0;	doodle_left_transparency_texture[49][48] = 0;	doodle_left_transparency_texture[49][49] = 0;	doodle_left_transparency_texture[49][50] = 0;	doodle_left_transparency_texture[49][51] = 0;	doodle_left_transparency_texture[49][52] = 0;	doodle_left_transparency_texture[49][53] = 0;	doodle_left_transparency_texture[49][54] = 0;	doodle_left_transparency_texture[49][55] = 0;	doodle_left_transparency_texture[49][56] = 0;	doodle_left_transparency_texture[49][57] = 0;	doodle_left_transparency_texture[49][58] = 0;	doodle_left_transparency_texture[49][59] = 0;	doodle_left_transparency_texture[49][60] = 0;	doodle_left_transparency_texture[49][61] = 0;	doodle_left_transparency_texture[49][62] = 0;	doodle_left_transparency_texture[49][63] = 0;	doodle_left_transparency_texture[49][64] = 0;	doodle_left_transparency_texture[49][65] = 0;	doodle_left_transparency_texture[49][66] = 0;	doodle_left_transparency_texture[49][67] = 0;	doodle_left_transparency_texture[49][68] = 0;	doodle_left_transparency_texture[49][69] = 0;	doodle_left_transparency_texture[49][70] = 0;	doodle_left_transparency_texture[49][71] = 0;	doodle_left_transparency_texture[49][72] = 0;	doodle_left_transparency_texture[49][73] = 0;	doodle_left_transparency_texture[49][74] = 0;	doodle_left_transparency_texture[49][75] = 0;	doodle_left_transparency_texture[49][76] = 1;	doodle_left_transparency_texture[49][77] = 1;	doodle_left_transparency_texture[49][78] = 1;	doodle_left_transparency_texture[49][79] = 1;	doodle_left_transparency_texture[50][0] = 1;	doodle_left_transparency_texture[50][1] = 1;	doodle_left_transparency_texture[50][2] = 1;	doodle_left_transparency_texture[50][3] = 1;	doodle_left_transparency_texture[50][4] = 1;	doodle_left_transparency_texture[50][5] = 1;	doodle_left_transparency_texture[50][6] = 1;	doodle_left_transparency_texture[50][7] = 1;	doodle_left_transparency_texture[50][8] = 1;	doodle_left_transparency_texture[50][9] = 1;	doodle_left_transparency_texture[50][10] = 1;	doodle_left_transparency_texture[50][11] = 1;	doodle_left_transparency_texture[50][12] = 1;	doodle_left_transparency_texture[50][13] = 1;	doodle_left_transparency_texture[50][14] = 1;	doodle_left_transparency_texture[50][15] = 1;	doodle_left_transparency_texture[50][16] = 1;	doodle_left_transparency_texture[50][17] = 1;	doodle_left_transparency_texture[50][18] = 1;	doodle_left_transparency_texture[50][19] = 1;	doodle_left_transparency_texture[50][20] = 1;	doodle_left_transparency_texture[50][21] = 1;	doodle_left_transparency_texture[50][22] = 1;	doodle_left_transparency_texture[50][23] = 1;	doodle_left_transparency_texture[50][24] = 1;	doodle_left_transparency_texture[50][25] = 1;	doodle_left_transparency_texture[50][26] = 1;	doodle_left_transparency_texture[50][27] = 1;	doodle_left_transparency_texture[50][28] = 0;	doodle_left_transparency_texture[50][29] = 0;	doodle_left_transparency_texture[50][30] = 0;	doodle_left_transparency_texture[50][31] = 0;	doodle_left_transparency_texture[50][32] = 0;	doodle_left_transparency_texture[50][33] = 0;	doodle_left_transparency_texture[50][34] = 0;	doodle_left_transparency_texture[50][35] = 0;	doodle_left_transparency_texture[50][36] = 0;	doodle_left_transparency_texture[50][37] = 0;	doodle_left_transparency_texture[50][38] = 0;	doodle_left_transparency_texture[50][39] = 0;	doodle_left_transparency_texture[50][40] = 0;	doodle_left_transparency_texture[50][41] = 0;	doodle_left_transparency_texture[50][42] = 0;	doodle_left_transparency_texture[50][43] = 0;	doodle_left_transparency_texture[50][44] = 0;	doodle_left_transparency_texture[50][45] = 0;	doodle_left_transparency_texture[50][46] = 0;	doodle_left_transparency_texture[50][47] = 0;	doodle_left_transparency_texture[50][48] = 0;	doodle_left_transparency_texture[50][49] = 0;	doodle_left_transparency_texture[50][50] = 0;	doodle_left_transparency_texture[50][51] = 0;	doodle_left_transparency_texture[50][52] = 0;	doodle_left_transparency_texture[50][53] = 0;	doodle_left_transparency_texture[50][54] = 0;	doodle_left_transparency_texture[50][55] = 0;	doodle_left_transparency_texture[50][56] = 0;	doodle_left_transparency_texture[50][57] = 0;	doodle_left_transparency_texture[50][58] = 0;	doodle_left_transparency_texture[50][59] = 0;	doodle_left_transparency_texture[50][60] = 0;	doodle_left_transparency_texture[50][61] = 0;	doodle_left_transparency_texture[50][62] = 0;	doodle_left_transparency_texture[50][63] = 0;	doodle_left_transparency_texture[50][64] = 0;	doodle_left_transparency_texture[50][65] = 0;	doodle_left_transparency_texture[50][66] = 0;	doodle_left_transparency_texture[50][67] = 0;	doodle_left_transparency_texture[50][68] = 0;	doodle_left_transparency_texture[50][69] = 0;	doodle_left_transparency_texture[50][70] = 0;	doodle_left_transparency_texture[50][71] = 0;	doodle_left_transparency_texture[50][72] = 0;	doodle_left_transparency_texture[50][73] = 0;	doodle_left_transparency_texture[50][74] = 0;	doodle_left_transparency_texture[50][75] = 0;	doodle_left_transparency_texture[50][76] = 1;	doodle_left_transparency_texture[50][77] = 1;	doodle_left_transparency_texture[50][78] = 1;	doodle_left_transparency_texture[50][79] = 1;	doodle_left_transparency_texture[51][0] = 1;	doodle_left_transparency_texture[51][1] = 1;	doodle_left_transparency_texture[51][2] = 1;	doodle_left_transparency_texture[51][3] = 1;	doodle_left_transparency_texture[51][4] = 1;	doodle_left_transparency_texture[51][5] = 1;	doodle_left_transparency_texture[51][6] = 1;	doodle_left_transparency_texture[51][7] = 1;	doodle_left_transparency_texture[51][8] = 1;	doodle_left_transparency_texture[51][9] = 1;	doodle_left_transparency_texture[51][10] = 1;	doodle_left_transparency_texture[51][11] = 1;	doodle_left_transparency_texture[51][12] = 1;	doodle_left_transparency_texture[51][13] = 1;	doodle_left_transparency_texture[51][14] = 1;	doodle_left_transparency_texture[51][15] = 1;	doodle_left_transparency_texture[51][16] = 1;	doodle_left_transparency_texture[51][17] = 1;	doodle_left_transparency_texture[51][18] = 1;	doodle_left_transparency_texture[51][19] = 1;	doodle_left_transparency_texture[51][20] = 1;	doodle_left_transparency_texture[51][21] = 1;	doodle_left_transparency_texture[51][22] = 1;	doodle_left_transparency_texture[51][23] = 1;	doodle_left_transparency_texture[51][24] = 1;	doodle_left_transparency_texture[51][25] = 1;	doodle_left_transparency_texture[51][26] = 1;	doodle_left_transparency_texture[51][27] = 1;	doodle_left_transparency_texture[51][28] = 0;	doodle_left_transparency_texture[51][29] = 0;	doodle_left_transparency_texture[51][30] = 0;	doodle_left_transparency_texture[51][31] = 0;	doodle_left_transparency_texture[51][32] = 0;	doodle_left_transparency_texture[51][33] = 0;	doodle_left_transparency_texture[51][34] = 0;	doodle_left_transparency_texture[51][35] = 0;	doodle_left_transparency_texture[51][36] = 0;	doodle_left_transparency_texture[51][37] = 0;	doodle_left_transparency_texture[51][38] = 0;	doodle_left_transparency_texture[51][39] = 0;	doodle_left_transparency_texture[51][40] = 0;	doodle_left_transparency_texture[51][41] = 0;	doodle_left_transparency_texture[51][42] = 0;	doodle_left_transparency_texture[51][43] = 0;	doodle_left_transparency_texture[51][44] = 0;	doodle_left_transparency_texture[51][45] = 0;	doodle_left_transparency_texture[51][46] = 0;	doodle_left_transparency_texture[51][47] = 0;	doodle_left_transparency_texture[51][48] = 0;	doodle_left_transparency_texture[51][49] = 0;	doodle_left_transparency_texture[51][50] = 0;	doodle_left_transparency_texture[51][51] = 0;	doodle_left_transparency_texture[51][52] = 0;	doodle_left_transparency_texture[51][53] = 0;	doodle_left_transparency_texture[51][54] = 0;	doodle_left_transparency_texture[51][55] = 0;	doodle_left_transparency_texture[51][56] = 0;	doodle_left_transparency_texture[51][57] = 0;	doodle_left_transparency_texture[51][58] = 0;	doodle_left_transparency_texture[51][59] = 0;	doodle_left_transparency_texture[51][60] = 0;	doodle_left_transparency_texture[51][61] = 0;	doodle_left_transparency_texture[51][62] = 0;	doodle_left_transparency_texture[51][63] = 0;	doodle_left_transparency_texture[51][64] = 0;	doodle_left_transparency_texture[51][65] = 0;	doodle_left_transparency_texture[51][66] = 0;	doodle_left_transparency_texture[51][67] = 0;	doodle_left_transparency_texture[51][68] = 0;	doodle_left_transparency_texture[51][69] = 0;	doodle_left_transparency_texture[51][70] = 0;	doodle_left_transparency_texture[51][71] = 0;	doodle_left_transparency_texture[51][72] = 0;	doodle_left_transparency_texture[51][73] = 0;	doodle_left_transparency_texture[51][74] = 0;	doodle_left_transparency_texture[51][75] = 0;	doodle_left_transparency_texture[51][76] = 1;	doodle_left_transparency_texture[51][77] = 1;	doodle_left_transparency_texture[51][78] = 1;	doodle_left_transparency_texture[51][79] = 1;	doodle_left_transparency_texture[52][0] = 1;	doodle_left_transparency_texture[52][1] = 1;	doodle_left_transparency_texture[52][2] = 1;	doodle_left_transparency_texture[52][3] = 1;	doodle_left_transparency_texture[52][4] = 1;	doodle_left_transparency_texture[52][5] = 1;	doodle_left_transparency_texture[52][6] = 1;	doodle_left_transparency_texture[52][7] = 1;	doodle_left_transparency_texture[52][8] = 1;	doodle_left_transparency_texture[52][9] = 1;	doodle_left_transparency_texture[52][10] = 1;	doodle_left_transparency_texture[52][11] = 1;	doodle_left_transparency_texture[52][12] = 1;	doodle_left_transparency_texture[52][13] = 1;	doodle_left_transparency_texture[52][14] = 1;	doodle_left_transparency_texture[52][15] = 1;	doodle_left_transparency_texture[52][16] = 1;	doodle_left_transparency_texture[52][17] = 1;	doodle_left_transparency_texture[52][18] = 1;	doodle_left_transparency_texture[52][19] = 1;	doodle_left_transparency_texture[52][20] = 1;	doodle_left_transparency_texture[52][21] = 1;	doodle_left_transparency_texture[52][22] = 1;	doodle_left_transparency_texture[52][23] = 1;	doodle_left_transparency_texture[52][24] = 1;	doodle_left_transparency_texture[52][25] = 1;	doodle_left_transparency_texture[52][26] = 1;	doodle_left_transparency_texture[52][27] = 1;	doodle_left_transparency_texture[52][28] = 0;	doodle_left_transparency_texture[52][29] = 0;	doodle_left_transparency_texture[52][30] = 0;	doodle_left_transparency_texture[52][31] = 0;	doodle_left_transparency_texture[52][32] = 0;	doodle_left_transparency_texture[52][33] = 0;	doodle_left_transparency_texture[52][34] = 0;	doodle_left_transparency_texture[52][35] = 0;	doodle_left_transparency_texture[52][36] = 0;	doodle_left_transparency_texture[52][37] = 0;	doodle_left_transparency_texture[52][38] = 0;	doodle_left_transparency_texture[52][39] = 0;	doodle_left_transparency_texture[52][40] = 0;	doodle_left_transparency_texture[52][41] = 0;	doodle_left_transparency_texture[52][42] = 0;	doodle_left_transparency_texture[52][43] = 0;	doodle_left_transparency_texture[52][44] = 0;	doodle_left_transparency_texture[52][45] = 0;	doodle_left_transparency_texture[52][46] = 0;	doodle_left_transparency_texture[52][47] = 0;	doodle_left_transparency_texture[52][48] = 0;	doodle_left_transparency_texture[52][49] = 0;	doodle_left_transparency_texture[52][50] = 0;	doodle_left_transparency_texture[52][51] = 0;	doodle_left_transparency_texture[52][52] = 0;	doodle_left_transparency_texture[52][53] = 0;	doodle_left_transparency_texture[52][54] = 0;	doodle_left_transparency_texture[52][55] = 0;	doodle_left_transparency_texture[52][56] = 0;	doodle_left_transparency_texture[52][57] = 0;	doodle_left_transparency_texture[52][58] = 0;	doodle_left_transparency_texture[52][59] = 0;	doodle_left_transparency_texture[52][60] = 0;	doodle_left_transparency_texture[52][61] = 0;	doodle_left_transparency_texture[52][62] = 0;	doodle_left_transparency_texture[52][63] = 0;	doodle_left_transparency_texture[52][64] = 0;	doodle_left_transparency_texture[52][65] = 0;	doodle_left_transparency_texture[52][66] = 0;	doodle_left_transparency_texture[52][67] = 0;	doodle_left_transparency_texture[52][68] = 0;	doodle_left_transparency_texture[52][69] = 0;	doodle_left_transparency_texture[52][70] = 0;	doodle_left_transparency_texture[52][71] = 0;	doodle_left_transparency_texture[52][72] = 0;	doodle_left_transparency_texture[52][73] = 0;	doodle_left_transparency_texture[52][74] = 0;	doodle_left_transparency_texture[52][75] = 0;	doodle_left_transparency_texture[52][76] = 1;	doodle_left_transparency_texture[52][77] = 1;	doodle_left_transparency_texture[52][78] = 1;	doodle_left_transparency_texture[52][79] = 1;	doodle_left_transparency_texture[53][0] = 1;	doodle_left_transparency_texture[53][1] = 1;	doodle_left_transparency_texture[53][2] = 1;	doodle_left_transparency_texture[53][3] = 1;	doodle_left_transparency_texture[53][4] = 1;	doodle_left_transparency_texture[53][5] = 1;	doodle_left_transparency_texture[53][6] = 1;	doodle_left_transparency_texture[53][7] = 1;	doodle_left_transparency_texture[53][8] = 1;	doodle_left_transparency_texture[53][9] = 1;	doodle_left_transparency_texture[53][10] = 1;	doodle_left_transparency_texture[53][11] = 1;	doodle_left_transparency_texture[53][12] = 1;	doodle_left_transparency_texture[53][13] = 1;	doodle_left_transparency_texture[53][14] = 1;	doodle_left_transparency_texture[53][15] = 1;	doodle_left_transparency_texture[53][16] = 1;	doodle_left_transparency_texture[53][17] = 1;	doodle_left_transparency_texture[53][18] = 1;	doodle_left_transparency_texture[53][19] = 1;	doodle_left_transparency_texture[53][20] = 1;	doodle_left_transparency_texture[53][21] = 1;	doodle_left_transparency_texture[53][22] = 1;	doodle_left_transparency_texture[53][23] = 1;	doodle_left_transparency_texture[53][24] = 1;	doodle_left_transparency_texture[53][25] = 1;	doodle_left_transparency_texture[53][26] = 1;	doodle_left_transparency_texture[53][27] = 1;	doodle_left_transparency_texture[53][28] = 0;	doodle_left_transparency_texture[53][29] = 0;	doodle_left_transparency_texture[53][30] = 0;	doodle_left_transparency_texture[53][31] = 0;	doodle_left_transparency_texture[53][32] = 0;	doodle_left_transparency_texture[53][33] = 0;	doodle_left_transparency_texture[53][34] = 0;	doodle_left_transparency_texture[53][35] = 0;	doodle_left_transparency_texture[53][36] = 0;	doodle_left_transparency_texture[53][37] = 0;	doodle_left_transparency_texture[53][38] = 0;	doodle_left_transparency_texture[53][39] = 0;	doodle_left_transparency_texture[53][40] = 0;	doodle_left_transparency_texture[53][41] = 0;	doodle_left_transparency_texture[53][42] = 0;	doodle_left_transparency_texture[53][43] = 0;	doodle_left_transparency_texture[53][44] = 0;	doodle_left_transparency_texture[53][45] = 0;	doodle_left_transparency_texture[53][46] = 0;	doodle_left_transparency_texture[53][47] = 0;	doodle_left_transparency_texture[53][48] = 0;	doodle_left_transparency_texture[53][49] = 0;	doodle_left_transparency_texture[53][50] = 0;	doodle_left_transparency_texture[53][51] = 0;	doodle_left_transparency_texture[53][52] = 0;	doodle_left_transparency_texture[53][53] = 0;	doodle_left_transparency_texture[53][54] = 0;	doodle_left_transparency_texture[53][55] = 0;	doodle_left_transparency_texture[53][56] = 0;	doodle_left_transparency_texture[53][57] = 0;	doodle_left_transparency_texture[53][58] = 0;	doodle_left_transparency_texture[53][59] = 0;	doodle_left_transparency_texture[53][60] = 0;	doodle_left_transparency_texture[53][61] = 0;	doodle_left_transparency_texture[53][62] = 0;	doodle_left_transparency_texture[53][63] = 0;	doodle_left_transparency_texture[53][64] = 0;	doodle_left_transparency_texture[53][65] = 0;	doodle_left_transparency_texture[53][66] = 0;	doodle_left_transparency_texture[53][67] = 0;	doodle_left_transparency_texture[53][68] = 0;	doodle_left_transparency_texture[53][69] = 0;	doodle_left_transparency_texture[53][70] = 0;	doodle_left_transparency_texture[53][71] = 0;	doodle_left_transparency_texture[53][72] = 0;	doodle_left_transparency_texture[53][73] = 0;	doodle_left_transparency_texture[53][74] = 0;	doodle_left_transparency_texture[53][75] = 0;	doodle_left_transparency_texture[53][76] = 1;	doodle_left_transparency_texture[53][77] = 1;	doodle_left_transparency_texture[53][78] = 1;	doodle_left_transparency_texture[53][79] = 1;	doodle_left_transparency_texture[54][0] = 1;	doodle_left_transparency_texture[54][1] = 1;	doodle_left_transparency_texture[54][2] = 1;	doodle_left_transparency_texture[54][3] = 1;	doodle_left_transparency_texture[54][4] = 1;	doodle_left_transparency_texture[54][5] = 1;	doodle_left_transparency_texture[54][6] = 1;	doodle_left_transparency_texture[54][7] = 1;	doodle_left_transparency_texture[54][8] = 1;	doodle_left_transparency_texture[54][9] = 1;	doodle_left_transparency_texture[54][10] = 1;	doodle_left_transparency_texture[54][11] = 1;	doodle_left_transparency_texture[54][12] = 1;	doodle_left_transparency_texture[54][13] = 1;	doodle_left_transparency_texture[54][14] = 1;	doodle_left_transparency_texture[54][15] = 1;	doodle_left_transparency_texture[54][16] = 1;	doodle_left_transparency_texture[54][17] = 1;	doodle_left_transparency_texture[54][18] = 1;	doodle_left_transparency_texture[54][19] = 1;	doodle_left_transparency_texture[54][20] = 1;	doodle_left_transparency_texture[54][21] = 1;	doodle_left_transparency_texture[54][22] = 1;	doodle_left_transparency_texture[54][23] = 1;	doodle_left_transparency_texture[54][24] = 1;	doodle_left_transparency_texture[54][25] = 1;	doodle_left_transparency_texture[54][26] = 1;	doodle_left_transparency_texture[54][27] = 1;	doodle_left_transparency_texture[54][28] = 0;	doodle_left_transparency_texture[54][29] = 0;	doodle_left_transparency_texture[54][30] = 0;	doodle_left_transparency_texture[54][31] = 0;	doodle_left_transparency_texture[54][32] = 0;	doodle_left_transparency_texture[54][33] = 0;	doodle_left_transparency_texture[54][34] = 0;	doodle_left_transparency_texture[54][35] = 0;	doodle_left_transparency_texture[54][36] = 0;	doodle_left_transparency_texture[54][37] = 0;	doodle_left_transparency_texture[54][38] = 0;	doodle_left_transparency_texture[54][39] = 0;	doodle_left_transparency_texture[54][40] = 0;	doodle_left_transparency_texture[54][41] = 0;	doodle_left_transparency_texture[54][42] = 0;	doodle_left_transparency_texture[54][43] = 0;	doodle_left_transparency_texture[54][44] = 0;	doodle_left_transparency_texture[54][45] = 0;	doodle_left_transparency_texture[54][46] = 0;	doodle_left_transparency_texture[54][47] = 0;	doodle_left_transparency_texture[54][48] = 0;	doodle_left_transparency_texture[54][49] = 0;	doodle_left_transparency_texture[54][50] = 0;	doodle_left_transparency_texture[54][51] = 0;	doodle_left_transparency_texture[54][52] = 0;	doodle_left_transparency_texture[54][53] = 0;	doodle_left_transparency_texture[54][54] = 0;	doodle_left_transparency_texture[54][55] = 0;	doodle_left_transparency_texture[54][56] = 0;	doodle_left_transparency_texture[54][57] = 0;	doodle_left_transparency_texture[54][58] = 0;	doodle_left_transparency_texture[54][59] = 0;	doodle_left_transparency_texture[54][60] = 0;	doodle_left_transparency_texture[54][61] = 0;	doodle_left_transparency_texture[54][62] = 0;	doodle_left_transparency_texture[54][63] = 0;	doodle_left_transparency_texture[54][64] = 0;	doodle_left_transparency_texture[54][65] = 0;	doodle_left_transparency_texture[54][66] = 0;	doodle_left_transparency_texture[54][67] = 0;	doodle_left_transparency_texture[54][68] = 0;	doodle_left_transparency_texture[54][69] = 0;	doodle_left_transparency_texture[54][70] = 0;	doodle_left_transparency_texture[54][71] = 0;	doodle_left_transparency_texture[54][72] = 0;	doodle_left_transparency_texture[54][73] = 0;	doodle_left_transparency_texture[54][74] = 0;	doodle_left_transparency_texture[54][75] = 0;	doodle_left_transparency_texture[54][76] = 1;	doodle_left_transparency_texture[54][77] = 1;	doodle_left_transparency_texture[54][78] = 1;	doodle_left_transparency_texture[54][79] = 1;	doodle_left_transparency_texture[55][0] = 1;	doodle_left_transparency_texture[55][1] = 1;	doodle_left_transparency_texture[55][2] = 1;	doodle_left_transparency_texture[55][3] = 1;	doodle_left_transparency_texture[55][4] = 1;	doodle_left_transparency_texture[55][5] = 1;	doodle_left_transparency_texture[55][6] = 1;	doodle_left_transparency_texture[55][7] = 1;	doodle_left_transparency_texture[55][8] = 1;	doodle_left_transparency_texture[55][9] = 1;	doodle_left_transparency_texture[55][10] = 1;	doodle_left_transparency_texture[55][11] = 1;	doodle_left_transparency_texture[55][12] = 1;	doodle_left_transparency_texture[55][13] = 1;	doodle_left_transparency_texture[55][14] = 1;	doodle_left_transparency_texture[55][15] = 1;	doodle_left_transparency_texture[55][16] = 1;	doodle_left_transparency_texture[55][17] = 1;	doodle_left_transparency_texture[55][18] = 1;	doodle_left_transparency_texture[55][19] = 1;	doodle_left_transparency_texture[55][20] = 1;	doodle_left_transparency_texture[55][21] = 1;	doodle_left_transparency_texture[55][22] = 1;	doodle_left_transparency_texture[55][23] = 1;	doodle_left_transparency_texture[55][24] = 1;	doodle_left_transparency_texture[55][25] = 1;	doodle_left_transparency_texture[55][26] = 1;	doodle_left_transparency_texture[55][27] = 1;	doodle_left_transparency_texture[55][28] = 0;	doodle_left_transparency_texture[55][29] = 0;	doodle_left_transparency_texture[55][30] = 0;	doodle_left_transparency_texture[55][31] = 0;	doodle_left_transparency_texture[55][32] = 0;	doodle_left_transparency_texture[55][33] = 0;	doodle_left_transparency_texture[55][34] = 0;	doodle_left_transparency_texture[55][35] = 0;	doodle_left_transparency_texture[55][36] = 0;	doodle_left_transparency_texture[55][37] = 0;	doodle_left_transparency_texture[55][38] = 0;	doodle_left_transparency_texture[55][39] = 0;	doodle_left_transparency_texture[55][40] = 0;	doodle_left_transparency_texture[55][41] = 0;	doodle_left_transparency_texture[55][42] = 0;	doodle_left_transparency_texture[55][43] = 0;	doodle_left_transparency_texture[55][44] = 0;	doodle_left_transparency_texture[55][45] = 0;	doodle_left_transparency_texture[55][46] = 0;	doodle_left_transparency_texture[55][47] = 0;	doodle_left_transparency_texture[55][48] = 0;	doodle_left_transparency_texture[55][49] = 0;	doodle_left_transparency_texture[55][50] = 0;	doodle_left_transparency_texture[55][51] = 0;	doodle_left_transparency_texture[55][52] = 0;	doodle_left_transparency_texture[55][53] = 0;	doodle_left_transparency_texture[55][54] = 0;	doodle_left_transparency_texture[55][55] = 0;	doodle_left_transparency_texture[55][56] = 0;	doodle_left_transparency_texture[55][57] = 0;	doodle_left_transparency_texture[55][58] = 0;	doodle_left_transparency_texture[55][59] = 0;	doodle_left_transparency_texture[55][60] = 0;	doodle_left_transparency_texture[55][61] = 0;	doodle_left_transparency_texture[55][62] = 0;	doodle_left_transparency_texture[55][63] = 0;	doodle_left_transparency_texture[55][64] = 0;	doodle_left_transparency_texture[55][65] = 0;	doodle_left_transparency_texture[55][66] = 0;	doodle_left_transparency_texture[55][67] = 0;	doodle_left_transparency_texture[55][68] = 0;	doodle_left_transparency_texture[55][69] = 0;	doodle_left_transparency_texture[55][70] = 0;	doodle_left_transparency_texture[55][71] = 0;	doodle_left_transparency_texture[55][72] = 0;	doodle_left_transparency_texture[55][73] = 0;	doodle_left_transparency_texture[55][74] = 0;	doodle_left_transparency_texture[55][75] = 0;	doodle_left_transparency_texture[55][76] = 1;	doodle_left_transparency_texture[55][77] = 1;	doodle_left_transparency_texture[55][78] = 1;	doodle_left_transparency_texture[55][79] = 1;	doodle_left_transparency_texture[56][0] = 1;	doodle_left_transparency_texture[56][1] = 1;	doodle_left_transparency_texture[56][2] = 1;	doodle_left_transparency_texture[56][3] = 1;	doodle_left_transparency_texture[56][4] = 1;	doodle_left_transparency_texture[56][5] = 1;	doodle_left_transparency_texture[56][6] = 1;	doodle_left_transparency_texture[56][7] = 1;	doodle_left_transparency_texture[56][8] = 1;	doodle_left_transparency_texture[56][9] = 1;	doodle_left_transparency_texture[56][10] = 1;	doodle_left_transparency_texture[56][11] = 1;	doodle_left_transparency_texture[56][12] = 1;	doodle_left_transparency_texture[56][13] = 1;	doodle_left_transparency_texture[56][14] = 1;	doodle_left_transparency_texture[56][15] = 1;	doodle_left_transparency_texture[56][16] = 1;	doodle_left_transparency_texture[56][17] = 1;	doodle_left_transparency_texture[56][18] = 1;	doodle_left_transparency_texture[56][19] = 1;	doodle_left_transparency_texture[56][20] = 1;	doodle_left_transparency_texture[56][21] = 1;	doodle_left_transparency_texture[56][22] = 1;	doodle_left_transparency_texture[56][23] = 1;	doodle_left_transparency_texture[56][24] = 1;	doodle_left_transparency_texture[56][25] = 1;	doodle_left_transparency_texture[56][26] = 1;	doodle_left_transparency_texture[56][27] = 1;	doodle_left_transparency_texture[56][28] = 0;	doodle_left_transparency_texture[56][29] = 0;	doodle_left_transparency_texture[56][30] = 0;	doodle_left_transparency_texture[56][31] = 0;	doodle_left_transparency_texture[56][32] = 0;	doodle_left_transparency_texture[56][33] = 0;	doodle_left_transparency_texture[56][34] = 0;	doodle_left_transparency_texture[56][35] = 0;	doodle_left_transparency_texture[56][36] = 0;	doodle_left_transparency_texture[56][37] = 0;	doodle_left_transparency_texture[56][38] = 0;	doodle_left_transparency_texture[56][39] = 0;	doodle_left_transparency_texture[56][40] = 0;	doodle_left_transparency_texture[56][41] = 0;	doodle_left_transparency_texture[56][42] = 0;	doodle_left_transparency_texture[56][43] = 0;	doodle_left_transparency_texture[56][44] = 0;	doodle_left_transparency_texture[56][45] = 0;	doodle_left_transparency_texture[56][46] = 0;	doodle_left_transparency_texture[56][47] = 0;	doodle_left_transparency_texture[56][48] = 0;	doodle_left_transparency_texture[56][49] = 0;	doodle_left_transparency_texture[56][50] = 0;	doodle_left_transparency_texture[56][51] = 0;	doodle_left_transparency_texture[56][52] = 0;	doodle_left_transparency_texture[56][53] = 0;	doodle_left_transparency_texture[56][54] = 0;	doodle_left_transparency_texture[56][55] = 0;	doodle_left_transparency_texture[56][56] = 0;	doodle_left_transparency_texture[56][57] = 0;	doodle_left_transparency_texture[56][58] = 0;	doodle_left_transparency_texture[56][59] = 0;	doodle_left_transparency_texture[56][60] = 0;	doodle_left_transparency_texture[56][61] = 0;	doodle_left_transparency_texture[56][62] = 0;	doodle_left_transparency_texture[56][63] = 0;	doodle_left_transparency_texture[56][64] = 0;	doodle_left_transparency_texture[56][65] = 0;	doodle_left_transparency_texture[56][66] = 0;	doodle_left_transparency_texture[56][67] = 0;	doodle_left_transparency_texture[56][68] = 0;	doodle_left_transparency_texture[56][69] = 0;	doodle_left_transparency_texture[56][70] = 0;	doodle_left_transparency_texture[56][71] = 0;	doodle_left_transparency_texture[56][72] = 0;	doodle_left_transparency_texture[56][73] = 0;	doodle_left_transparency_texture[56][74] = 0;	doodle_left_transparency_texture[56][75] = 0;	doodle_left_transparency_texture[56][76] = 1;	doodle_left_transparency_texture[56][77] = 1;	doodle_left_transparency_texture[56][78] = 1;	doodle_left_transparency_texture[56][79] = 1;	doodle_left_transparency_texture[57][0] = 1;	doodle_left_transparency_texture[57][1] = 1;	doodle_left_transparency_texture[57][2] = 1;	doodle_left_transparency_texture[57][3] = 1;	doodle_left_transparency_texture[57][4] = 1;	doodle_left_transparency_texture[57][5] = 1;	doodle_left_transparency_texture[57][6] = 1;	doodle_left_transparency_texture[57][7] = 1;	doodle_left_transparency_texture[57][8] = 1;	doodle_left_transparency_texture[57][9] = 1;	doodle_left_transparency_texture[57][10] = 1;	doodle_left_transparency_texture[57][11] = 1;	doodle_left_transparency_texture[57][12] = 1;	doodle_left_transparency_texture[57][13] = 1;	doodle_left_transparency_texture[57][14] = 1;	doodle_left_transparency_texture[57][15] = 1;	doodle_left_transparency_texture[57][16] = 1;	doodle_left_transparency_texture[57][17] = 1;	doodle_left_transparency_texture[57][18] = 1;	doodle_left_transparency_texture[57][19] = 1;	doodle_left_transparency_texture[57][20] = 1;	doodle_left_transparency_texture[57][21] = 1;	doodle_left_transparency_texture[57][22] = 1;	doodle_left_transparency_texture[57][23] = 1;	doodle_left_transparency_texture[57][24] = 1;	doodle_left_transparency_texture[57][25] = 1;	doodle_left_transparency_texture[57][26] = 1;	doodle_left_transparency_texture[57][27] = 1;	doodle_left_transparency_texture[57][28] = 0;	doodle_left_transparency_texture[57][29] = 0;	doodle_left_transparency_texture[57][30] = 0;	doodle_left_transparency_texture[57][31] = 0;	doodle_left_transparency_texture[57][32] = 0;	doodle_left_transparency_texture[57][33] = 0;	doodle_left_transparency_texture[57][34] = 0;	doodle_left_transparency_texture[57][35] = 0;	doodle_left_transparency_texture[57][36] = 0;	doodle_left_transparency_texture[57][37] = 0;	doodle_left_transparency_texture[57][38] = 0;	doodle_left_transparency_texture[57][39] = 0;	doodle_left_transparency_texture[57][40] = 0;	doodle_left_transparency_texture[57][41] = 0;	doodle_left_transparency_texture[57][42] = 0;	doodle_left_transparency_texture[57][43] = 0;	doodle_left_transparency_texture[57][44] = 0;	doodle_left_transparency_texture[57][45] = 0;	doodle_left_transparency_texture[57][46] = 0;	doodle_left_transparency_texture[57][47] = 0;	doodle_left_transparency_texture[57][48] = 0;	doodle_left_transparency_texture[57][49] = 0;	doodle_left_transparency_texture[57][50] = 0;	doodle_left_transparency_texture[57][51] = 0;	doodle_left_transparency_texture[57][52] = 0;	doodle_left_transparency_texture[57][53] = 0;	doodle_left_transparency_texture[57][54] = 0;	doodle_left_transparency_texture[57][55] = 0;	doodle_left_transparency_texture[57][56] = 0;	doodle_left_transparency_texture[57][57] = 0;	doodle_left_transparency_texture[57][58] = 0;	doodle_left_transparency_texture[57][59] = 0;	doodle_left_transparency_texture[57][60] = 0;	doodle_left_transparency_texture[57][61] = 0;	doodle_left_transparency_texture[57][62] = 0;	doodle_left_transparency_texture[57][63] = 0;	doodle_left_transparency_texture[57][64] = 0;	doodle_left_transparency_texture[57][65] = 0;	doodle_left_transparency_texture[57][66] = 0;	doodle_left_transparency_texture[57][67] = 0;	doodle_left_transparency_texture[57][68] = 0;	doodle_left_transparency_texture[57][69] = 0;	doodle_left_transparency_texture[57][70] = 0;	doodle_left_transparency_texture[57][71] = 0;	doodle_left_transparency_texture[57][72] = 0;	doodle_left_transparency_texture[57][73] = 0;	doodle_left_transparency_texture[57][74] = 0;	doodle_left_transparency_texture[57][75] = 0;	doodle_left_transparency_texture[57][76] = 1;	doodle_left_transparency_texture[57][77] = 1;	doodle_left_transparency_texture[57][78] = 1;	doodle_left_transparency_texture[57][79] = 1;	doodle_left_transparency_texture[58][0] = 1;	doodle_left_transparency_texture[58][1] = 1;	doodle_left_transparency_texture[58][2] = 1;	doodle_left_transparency_texture[58][3] = 1;	doodle_left_transparency_texture[58][4] = 1;	doodle_left_transparency_texture[58][5] = 1;	doodle_left_transparency_texture[58][6] = 1;	doodle_left_transparency_texture[58][7] = 1;	doodle_left_transparency_texture[58][8] = 1;	doodle_left_transparency_texture[58][9] = 1;	doodle_left_transparency_texture[58][10] = 1;	doodle_left_transparency_texture[58][11] = 1;	doodle_left_transparency_texture[58][12] = 1;	doodle_left_transparency_texture[58][13] = 1;	doodle_left_transparency_texture[58][14] = 1;	doodle_left_transparency_texture[58][15] = 1;	doodle_left_transparency_texture[58][16] = 1;	doodle_left_transparency_texture[58][17] = 1;	doodle_left_transparency_texture[58][18] = 1;	doodle_left_transparency_texture[58][19] = 1;	doodle_left_transparency_texture[58][20] = 1;	doodle_left_transparency_texture[58][21] = 1;	doodle_left_transparency_texture[58][22] = 1;	doodle_left_transparency_texture[58][23] = 1;	doodle_left_transparency_texture[58][24] = 1;	doodle_left_transparency_texture[58][25] = 1;	doodle_left_transparency_texture[58][26] = 1;	doodle_left_transparency_texture[58][27] = 1;	doodle_left_transparency_texture[58][28] = 0;	doodle_left_transparency_texture[58][29] = 0;	doodle_left_transparency_texture[58][30] = 0;	doodle_left_transparency_texture[58][31] = 0;	doodle_left_transparency_texture[58][32] = 0;	doodle_left_transparency_texture[58][33] = 0;	doodle_left_transparency_texture[58][34] = 0;	doodle_left_transparency_texture[58][35] = 0;	doodle_left_transparency_texture[58][36] = 0;	doodle_left_transparency_texture[58][37] = 0;	doodle_left_transparency_texture[58][38] = 0;	doodle_left_transparency_texture[58][39] = 0;	doodle_left_transparency_texture[58][40] = 0;	doodle_left_transparency_texture[58][41] = 0;	doodle_left_transparency_texture[58][42] = 0;	doodle_left_transparency_texture[58][43] = 0;	doodle_left_transparency_texture[58][44] = 0;	doodle_left_transparency_texture[58][45] = 0;	doodle_left_transparency_texture[58][46] = 0;	doodle_left_transparency_texture[58][47] = 0;	doodle_left_transparency_texture[58][48] = 0;	doodle_left_transparency_texture[58][49] = 0;	doodle_left_transparency_texture[58][50] = 0;	doodle_left_transparency_texture[58][51] = 0;	doodle_left_transparency_texture[58][52] = 0;	doodle_left_transparency_texture[58][53] = 0;	doodle_left_transparency_texture[58][54] = 0;	doodle_left_transparency_texture[58][55] = 0;	doodle_left_transparency_texture[58][56] = 0;	doodle_left_transparency_texture[58][57] = 0;	doodle_left_transparency_texture[58][58] = 0;	doodle_left_transparency_texture[58][59] = 0;	doodle_left_transparency_texture[58][60] = 0;	doodle_left_transparency_texture[58][61] = 0;	doodle_left_transparency_texture[58][62] = 0;	doodle_left_transparency_texture[58][63] = 0;	doodle_left_transparency_texture[58][64] = 0;	doodle_left_transparency_texture[58][65] = 0;	doodle_left_transparency_texture[58][66] = 0;	doodle_left_transparency_texture[58][67] = 0;	doodle_left_transparency_texture[58][68] = 0;	doodle_left_transparency_texture[58][69] = 0;	doodle_left_transparency_texture[58][70] = 0;	doodle_left_transparency_texture[58][71] = 0;	doodle_left_transparency_texture[58][72] = 0;	doodle_left_transparency_texture[58][73] = 0;	doodle_left_transparency_texture[58][74] = 0;	doodle_left_transparency_texture[58][75] = 0;	doodle_left_transparency_texture[58][76] = 1;	doodle_left_transparency_texture[58][77] = 1;	doodle_left_transparency_texture[58][78] = 1;	doodle_left_transparency_texture[58][79] = 1;	doodle_left_transparency_texture[59][0] = 1;	doodle_left_transparency_texture[59][1] = 1;	doodle_left_transparency_texture[59][2] = 1;	doodle_left_transparency_texture[59][3] = 1;	doodle_left_transparency_texture[59][4] = 1;	doodle_left_transparency_texture[59][5] = 1;	doodle_left_transparency_texture[59][6] = 1;	doodle_left_transparency_texture[59][7] = 1;	doodle_left_transparency_texture[59][8] = 1;	doodle_left_transparency_texture[59][9] = 1;	doodle_left_transparency_texture[59][10] = 1;	doodle_left_transparency_texture[59][11] = 1;	doodle_left_transparency_texture[59][12] = 1;	doodle_left_transparency_texture[59][13] = 1;	doodle_left_transparency_texture[59][14] = 1;	doodle_left_transparency_texture[59][15] = 1;	doodle_left_transparency_texture[59][16] = 1;	doodle_left_transparency_texture[59][17] = 1;	doodle_left_transparency_texture[59][18] = 1;	doodle_left_transparency_texture[59][19] = 1;	doodle_left_transparency_texture[59][20] = 1;	doodle_left_transparency_texture[59][21] = 1;	doodle_left_transparency_texture[59][22] = 1;	doodle_left_transparency_texture[59][23] = 1;	doodle_left_transparency_texture[59][24] = 1;	doodle_left_transparency_texture[59][25] = 1;	doodle_left_transparency_texture[59][26] = 1;	doodle_left_transparency_texture[59][27] = 1;	doodle_left_transparency_texture[59][28] = 0;	doodle_left_transparency_texture[59][29] = 0;	doodle_left_transparency_texture[59][30] = 0;	doodle_left_transparency_texture[59][31] = 0;	doodle_left_transparency_texture[59][32] = 0;	doodle_left_transparency_texture[59][33] = 0;	doodle_left_transparency_texture[59][34] = 0;	doodle_left_transparency_texture[59][35] = 0;	doodle_left_transparency_texture[59][36] = 0;	doodle_left_transparency_texture[59][37] = 0;	doodle_left_transparency_texture[59][38] = 0;	doodle_left_transparency_texture[59][39] = 0;	doodle_left_transparency_texture[59][40] = 0;	doodle_left_transparency_texture[59][41] = 0;	doodle_left_transparency_texture[59][42] = 0;	doodle_left_transparency_texture[59][43] = 0;	doodle_left_transparency_texture[59][44] = 0;	doodle_left_transparency_texture[59][45] = 0;	doodle_left_transparency_texture[59][46] = 0;	doodle_left_transparency_texture[59][47] = 0;	doodle_left_transparency_texture[59][48] = 0;	doodle_left_transparency_texture[59][49] = 0;	doodle_left_transparency_texture[59][50] = 0;	doodle_left_transparency_texture[59][51] = 0;	doodle_left_transparency_texture[59][52] = 0;	doodle_left_transparency_texture[59][53] = 0;	doodle_left_transparency_texture[59][54] = 0;	doodle_left_transparency_texture[59][55] = 0;	doodle_left_transparency_texture[59][56] = 0;	doodle_left_transparency_texture[59][57] = 0;	doodle_left_transparency_texture[59][58] = 0;	doodle_left_transparency_texture[59][59] = 0;	doodle_left_transparency_texture[59][60] = 0;	doodle_left_transparency_texture[59][61] = 0;	doodle_left_transparency_texture[59][62] = 0;	doodle_left_transparency_texture[59][63] = 0;	doodle_left_transparency_texture[59][64] = 0;	doodle_left_transparency_texture[59][65] = 0;	doodle_left_transparency_texture[59][66] = 0;	doodle_left_transparency_texture[59][67] = 0;	doodle_left_transparency_texture[59][68] = 0;	doodle_left_transparency_texture[59][69] = 0;	doodle_left_transparency_texture[59][70] = 0;	doodle_left_transparency_texture[59][71] = 0;	doodle_left_transparency_texture[59][72] = 0;	doodle_left_transparency_texture[59][73] = 0;	doodle_left_transparency_texture[59][74] = 0;	doodle_left_transparency_texture[59][75] = 0;	doodle_left_transparency_texture[59][76] = 1;	doodle_left_transparency_texture[59][77] = 1;	doodle_left_transparency_texture[59][78] = 1;	doodle_left_transparency_texture[59][79] = 1;	doodle_left_transparency_texture[60][0] = 1;	doodle_left_transparency_texture[60][1] = 1;	doodle_left_transparency_texture[60][2] = 1;	doodle_left_transparency_texture[60][3] = 1;	doodle_left_transparency_texture[60][4] = 1;	doodle_left_transparency_texture[60][5] = 1;	doodle_left_transparency_texture[60][6] = 1;	doodle_left_transparency_texture[60][7] = 1;	doodle_left_transparency_texture[60][8] = 1;	doodle_left_transparency_texture[60][9] = 1;	doodle_left_transparency_texture[60][10] = 1;	doodle_left_transparency_texture[60][11] = 1;	doodle_left_transparency_texture[60][12] = 1;	doodle_left_transparency_texture[60][13] = 1;	doodle_left_transparency_texture[60][14] = 1;	doodle_left_transparency_texture[60][15] = 1;	doodle_left_transparency_texture[60][16] = 1;	doodle_left_transparency_texture[60][17] = 1;	doodle_left_transparency_texture[60][18] = 1;	doodle_left_transparency_texture[60][19] = 1;	doodle_left_transparency_texture[60][20] = 1;	doodle_left_transparency_texture[60][21] = 1;	doodle_left_transparency_texture[60][22] = 1;	doodle_left_transparency_texture[60][23] = 1;	doodle_left_transparency_texture[60][24] = 1;	doodle_left_transparency_texture[60][25] = 1;	doodle_left_transparency_texture[60][26] = 1;	doodle_left_transparency_texture[60][27] = 1;	doodle_left_transparency_texture[60][28] = 1;	doodle_left_transparency_texture[60][29] = 1;	doodle_left_transparency_texture[60][30] = 1;	doodle_left_transparency_texture[60][31] = 1;	doodle_left_transparency_texture[60][32] = 0;	doodle_left_transparency_texture[60][33] = 0;	doodle_left_transparency_texture[60][34] = 0;	doodle_left_transparency_texture[60][35] = 0;	doodle_left_transparency_texture[60][36] = 1;	doodle_left_transparency_texture[60][37] = 1;	doodle_left_transparency_texture[60][38] = 1;	doodle_left_transparency_texture[60][39] = 1;	doodle_left_transparency_texture[60][40] = 1;	doodle_left_transparency_texture[60][41] = 1;	doodle_left_transparency_texture[60][42] = 1;	doodle_left_transparency_texture[60][43] = 1;	doodle_left_transparency_texture[60][44] = 0;	doodle_left_transparency_texture[60][45] = 0;	doodle_left_transparency_texture[60][46] = 0;	doodle_left_transparency_texture[60][47] = 0;	doodle_left_transparency_texture[60][48] = 1;	doodle_left_transparency_texture[60][49] = 1;	doodle_left_transparency_texture[60][50] = 1;	doodle_left_transparency_texture[60][51] = 1;	doodle_left_transparency_texture[60][52] = 1;	doodle_left_transparency_texture[60][53] = 1;	doodle_left_transparency_texture[60][54] = 1;	doodle_left_transparency_texture[60][55] = 1;	doodle_left_transparency_texture[60][56] = 0;	doodle_left_transparency_texture[60][57] = 0;	doodle_left_transparency_texture[60][58] = 0;	doodle_left_transparency_texture[60][59] = 0;	doodle_left_transparency_texture[60][60] = 1;	doodle_left_transparency_texture[60][61] = 1;	doodle_left_transparency_texture[60][62] = 1;	doodle_left_transparency_texture[60][63] = 1;	doodle_left_transparency_texture[60][64] = 1;	doodle_left_transparency_texture[60][65] = 1;	doodle_left_transparency_texture[60][66] = 1;	doodle_left_transparency_texture[60][67] = 1;	doodle_left_transparency_texture[60][68] = 0;	doodle_left_transparency_texture[60][69] = 0;	doodle_left_transparency_texture[60][70] = 0;	doodle_left_transparency_texture[60][71] = 0;	doodle_left_transparency_texture[60][72] = 1;	doodle_left_transparency_texture[60][73] = 1;	doodle_left_transparency_texture[60][74] = 1;	doodle_left_transparency_texture[60][75] = 1;	doodle_left_transparency_texture[60][76] = 1;	doodle_left_transparency_texture[60][77] = 1;	doodle_left_transparency_texture[60][78] = 1;	doodle_left_transparency_texture[60][79] = 1;	doodle_left_transparency_texture[61][0] = 1;	doodle_left_transparency_texture[61][1] = 1;	doodle_left_transparency_texture[61][2] = 1;	doodle_left_transparency_texture[61][3] = 1;	doodle_left_transparency_texture[61][4] = 1;	doodle_left_transparency_texture[61][5] = 1;	doodle_left_transparency_texture[61][6] = 1;	doodle_left_transparency_texture[61][7] = 1;	doodle_left_transparency_texture[61][8] = 1;	doodle_left_transparency_texture[61][9] = 1;	doodle_left_transparency_texture[61][10] = 1;	doodle_left_transparency_texture[61][11] = 1;	doodle_left_transparency_texture[61][12] = 1;	doodle_left_transparency_texture[61][13] = 1;	doodle_left_transparency_texture[61][14] = 1;	doodle_left_transparency_texture[61][15] = 1;	doodle_left_transparency_texture[61][16] = 1;	doodle_left_transparency_texture[61][17] = 1;	doodle_left_transparency_texture[61][18] = 1;	doodle_left_transparency_texture[61][19] = 1;	doodle_left_transparency_texture[61][20] = 1;	doodle_left_transparency_texture[61][21] = 1;	doodle_left_transparency_texture[61][22] = 1;	doodle_left_transparency_texture[61][23] = 1;	doodle_left_transparency_texture[61][24] = 1;	doodle_left_transparency_texture[61][25] = 1;	doodle_left_transparency_texture[61][26] = 1;	doodle_left_transparency_texture[61][27] = 1;	doodle_left_transparency_texture[61][28] = 1;	doodle_left_transparency_texture[61][29] = 1;	doodle_left_transparency_texture[61][30] = 1;	doodle_left_transparency_texture[61][31] = 1;	doodle_left_transparency_texture[61][32] = 0;	doodle_left_transparency_texture[61][33] = 0;	doodle_left_transparency_texture[61][34] = 0;	doodle_left_transparency_texture[61][35] = 0;	doodle_left_transparency_texture[61][36] = 1;	doodle_left_transparency_texture[61][37] = 1;	doodle_left_transparency_texture[61][38] = 1;	doodle_left_transparency_texture[61][39] = 1;	doodle_left_transparency_texture[61][40] = 1;	doodle_left_transparency_texture[61][41] = 1;	doodle_left_transparency_texture[61][42] = 1;	doodle_left_transparency_texture[61][43] = 1;	doodle_left_transparency_texture[61][44] = 0;	doodle_left_transparency_texture[61][45] = 0;	doodle_left_transparency_texture[61][46] = 0;	doodle_left_transparency_texture[61][47] = 0;	doodle_left_transparency_texture[61][48] = 1;	doodle_left_transparency_texture[61][49] = 1;	doodle_left_transparency_texture[61][50] = 1;	doodle_left_transparency_texture[61][51] = 1;	doodle_left_transparency_texture[61][52] = 1;	doodle_left_transparency_texture[61][53] = 1;	doodle_left_transparency_texture[61][54] = 1;	doodle_left_transparency_texture[61][55] = 1;	doodle_left_transparency_texture[61][56] = 0;	doodle_left_transparency_texture[61][57] = 0;	doodle_left_transparency_texture[61][58] = 0;	doodle_left_transparency_texture[61][59] = 0;	doodle_left_transparency_texture[61][60] = 1;	doodle_left_transparency_texture[61][61] = 1;	doodle_left_transparency_texture[61][62] = 1;	doodle_left_transparency_texture[61][63] = 1;	doodle_left_transparency_texture[61][64] = 1;	doodle_left_transparency_texture[61][65] = 1;	doodle_left_transparency_texture[61][66] = 1;	doodle_left_transparency_texture[61][67] = 1;	doodle_left_transparency_texture[61][68] = 0;	doodle_left_transparency_texture[61][69] = 0;	doodle_left_transparency_texture[61][70] = 0;	doodle_left_transparency_texture[61][71] = 0;	doodle_left_transparency_texture[61][72] = 1;	doodle_left_transparency_texture[61][73] = 1;	doodle_left_transparency_texture[61][74] = 1;	doodle_left_transparency_texture[61][75] = 1;	doodle_left_transparency_texture[61][76] = 1;	doodle_left_transparency_texture[61][77] = 1;	doodle_left_transparency_texture[61][78] = 1;	doodle_left_transparency_texture[61][79] = 1;	doodle_left_transparency_texture[62][0] = 1;	doodle_left_transparency_texture[62][1] = 1;	doodle_left_transparency_texture[62][2] = 1;	doodle_left_transparency_texture[62][3] = 1;	doodle_left_transparency_texture[62][4] = 1;	doodle_left_transparency_texture[62][5] = 1;	doodle_left_transparency_texture[62][6] = 1;	doodle_left_transparency_texture[62][7] = 1;	doodle_left_transparency_texture[62][8] = 1;	doodle_left_transparency_texture[62][9] = 1;	doodle_left_transparency_texture[62][10] = 1;	doodle_left_transparency_texture[62][11] = 1;	doodle_left_transparency_texture[62][12] = 1;	doodle_left_transparency_texture[62][13] = 1;	doodle_left_transparency_texture[62][14] = 1;	doodle_left_transparency_texture[62][15] = 1;	doodle_left_transparency_texture[62][16] = 1;	doodle_left_transparency_texture[62][17] = 1;	doodle_left_transparency_texture[62][18] = 1;	doodle_left_transparency_texture[62][19] = 1;	doodle_left_transparency_texture[62][20] = 1;	doodle_left_transparency_texture[62][21] = 1;	doodle_left_transparency_texture[62][22] = 1;	doodle_left_transparency_texture[62][23] = 1;	doodle_left_transparency_texture[62][24] = 1;	doodle_left_transparency_texture[62][25] = 1;	doodle_left_transparency_texture[62][26] = 1;	doodle_left_transparency_texture[62][27] = 1;	doodle_left_transparency_texture[62][28] = 1;	doodle_left_transparency_texture[62][29] = 1;	doodle_left_transparency_texture[62][30] = 1;	doodle_left_transparency_texture[62][31] = 1;	doodle_left_transparency_texture[62][32] = 0;	doodle_left_transparency_texture[62][33] = 0;	doodle_left_transparency_texture[62][34] = 0;	doodle_left_transparency_texture[62][35] = 0;	doodle_left_transparency_texture[62][36] = 1;	doodle_left_transparency_texture[62][37] = 1;	doodle_left_transparency_texture[62][38] = 1;	doodle_left_transparency_texture[62][39] = 1;	doodle_left_transparency_texture[62][40] = 1;	doodle_left_transparency_texture[62][41] = 1;	doodle_left_transparency_texture[62][42] = 1;	doodle_left_transparency_texture[62][43] = 1;	doodle_left_transparency_texture[62][44] = 0;	doodle_left_transparency_texture[62][45] = 0;	doodle_left_transparency_texture[62][46] = 0;	doodle_left_transparency_texture[62][47] = 0;	doodle_left_transparency_texture[62][48] = 1;	doodle_left_transparency_texture[62][49] = 1;	doodle_left_transparency_texture[62][50] = 1;	doodle_left_transparency_texture[62][51] = 1;	doodle_left_transparency_texture[62][52] = 1;	doodle_left_transparency_texture[62][53] = 1;	doodle_left_transparency_texture[62][54] = 1;	doodle_left_transparency_texture[62][55] = 1;	doodle_left_transparency_texture[62][56] = 0;	doodle_left_transparency_texture[62][57] = 0;	doodle_left_transparency_texture[62][58] = 0;	doodle_left_transparency_texture[62][59] = 0;	doodle_left_transparency_texture[62][60] = 1;	doodle_left_transparency_texture[62][61] = 1;	doodle_left_transparency_texture[62][62] = 1;	doodle_left_transparency_texture[62][63] = 1;	doodle_left_transparency_texture[62][64] = 1;	doodle_left_transparency_texture[62][65] = 1;	doodle_left_transparency_texture[62][66] = 1;	doodle_left_transparency_texture[62][67] = 1;	doodle_left_transparency_texture[62][68] = 0;	doodle_left_transparency_texture[62][69] = 0;	doodle_left_transparency_texture[62][70] = 0;	doodle_left_transparency_texture[62][71] = 0;	doodle_left_transparency_texture[62][72] = 1;	doodle_left_transparency_texture[62][73] = 1;	doodle_left_transparency_texture[62][74] = 1;	doodle_left_transparency_texture[62][75] = 1;	doodle_left_transparency_texture[62][76] = 1;	doodle_left_transparency_texture[62][77] = 1;	doodle_left_transparency_texture[62][78] = 1;	doodle_left_transparency_texture[62][79] = 1;	doodle_left_transparency_texture[63][0] = 1;	doodle_left_transparency_texture[63][1] = 1;	doodle_left_transparency_texture[63][2] = 1;	doodle_left_transparency_texture[63][3] = 1;	doodle_left_transparency_texture[63][4] = 1;	doodle_left_transparency_texture[63][5] = 1;	doodle_left_transparency_texture[63][6] = 1;	doodle_left_transparency_texture[63][7] = 1;	doodle_left_transparency_texture[63][8] = 1;	doodle_left_transparency_texture[63][9] = 1;	doodle_left_transparency_texture[63][10] = 1;	doodle_left_transparency_texture[63][11] = 1;	doodle_left_transparency_texture[63][12] = 1;	doodle_left_transparency_texture[63][13] = 1;	doodle_left_transparency_texture[63][14] = 1;	doodle_left_transparency_texture[63][15] = 1;	doodle_left_transparency_texture[63][16] = 1;	doodle_left_transparency_texture[63][17] = 1;	doodle_left_transparency_texture[63][18] = 1;	doodle_left_transparency_texture[63][19] = 1;	doodle_left_transparency_texture[63][20] = 1;	doodle_left_transparency_texture[63][21] = 1;	doodle_left_transparency_texture[63][22] = 1;	doodle_left_transparency_texture[63][23] = 1;	doodle_left_transparency_texture[63][24] = 1;	doodle_left_transparency_texture[63][25] = 1;	doodle_left_transparency_texture[63][26] = 1;	doodle_left_transparency_texture[63][27] = 1;	doodle_left_transparency_texture[63][28] = 1;	doodle_left_transparency_texture[63][29] = 1;	doodle_left_transparency_texture[63][30] = 1;	doodle_left_transparency_texture[63][31] = 1;	doodle_left_transparency_texture[63][32] = 0;	doodle_left_transparency_texture[63][33] = 0;	doodle_left_transparency_texture[63][34] = 0;	doodle_left_transparency_texture[63][35] = 0;	doodle_left_transparency_texture[63][36] = 1;	doodle_left_transparency_texture[63][37] = 1;	doodle_left_transparency_texture[63][38] = 1;	doodle_left_transparency_texture[63][39] = 1;	doodle_left_transparency_texture[63][40] = 1;	doodle_left_transparency_texture[63][41] = 1;	doodle_left_transparency_texture[63][42] = 1;	doodle_left_transparency_texture[63][43] = 1;	doodle_left_transparency_texture[63][44] = 0;	doodle_left_transparency_texture[63][45] = 0;	doodle_left_transparency_texture[63][46] = 0;	doodle_left_transparency_texture[63][47] = 0;	doodle_left_transparency_texture[63][48] = 1;	doodle_left_transparency_texture[63][49] = 1;	doodle_left_transparency_texture[63][50] = 1;	doodle_left_transparency_texture[63][51] = 1;	doodle_left_transparency_texture[63][52] = 1;	doodle_left_transparency_texture[63][53] = 1;	doodle_left_transparency_texture[63][54] = 1;	doodle_left_transparency_texture[63][55] = 1;	doodle_left_transparency_texture[63][56] = 0;	doodle_left_transparency_texture[63][57] = 0;	doodle_left_transparency_texture[63][58] = 0;	doodle_left_transparency_texture[63][59] = 0;	doodle_left_transparency_texture[63][60] = 1;	doodle_left_transparency_texture[63][61] = 1;	doodle_left_transparency_texture[63][62] = 1;	doodle_left_transparency_texture[63][63] = 1;	doodle_left_transparency_texture[63][64] = 1;	doodle_left_transparency_texture[63][65] = 1;	doodle_left_transparency_texture[63][66] = 1;	doodle_left_transparency_texture[63][67] = 1;	doodle_left_transparency_texture[63][68] = 0;	doodle_left_transparency_texture[63][69] = 0;	doodle_left_transparency_texture[63][70] = 0;	doodle_left_transparency_texture[63][71] = 0;	doodle_left_transparency_texture[63][72] = 1;	doodle_left_transparency_texture[63][73] = 1;	doodle_left_transparency_texture[63][74] = 1;	doodle_left_transparency_texture[63][75] = 1;	doodle_left_transparency_texture[63][76] = 1;	doodle_left_transparency_texture[63][77] = 1;	doodle_left_transparency_texture[63][78] = 1;	doodle_left_transparency_texture[63][79] = 1;	doodle_left_transparency_texture[64][0] = 1;	doodle_left_transparency_texture[64][1] = 1;	doodle_left_transparency_texture[64][2] = 1;	doodle_left_transparency_texture[64][3] = 1;	doodle_left_transparency_texture[64][4] = 1;	doodle_left_transparency_texture[64][5] = 1;	doodle_left_transparency_texture[64][6] = 1;	doodle_left_transparency_texture[64][7] = 1;	doodle_left_transparency_texture[64][8] = 1;	doodle_left_transparency_texture[64][9] = 1;	doodle_left_transparency_texture[64][10] = 1;	doodle_left_transparency_texture[64][11] = 1;	doodle_left_transparency_texture[64][12] = 1;	doodle_left_transparency_texture[64][13] = 1;	doodle_left_transparency_texture[64][14] = 1;	doodle_left_transparency_texture[64][15] = 1;	doodle_left_transparency_texture[64][16] = 1;	doodle_left_transparency_texture[64][17] = 1;	doodle_left_transparency_texture[64][18] = 1;	doodle_left_transparency_texture[64][19] = 1;	doodle_left_transparency_texture[64][20] = 1;	doodle_left_transparency_texture[64][21] = 1;	doodle_left_transparency_texture[64][22] = 1;	doodle_left_transparency_texture[64][23] = 1;	doodle_left_transparency_texture[64][24] = 1;	doodle_left_transparency_texture[64][25] = 1;	doodle_left_transparency_texture[64][26] = 1;	doodle_left_transparency_texture[64][27] = 1;	doodle_left_transparency_texture[64][28] = 1;	doodle_left_transparency_texture[64][29] = 1;	doodle_left_transparency_texture[64][30] = 1;	doodle_left_transparency_texture[64][31] = 1;	doodle_left_transparency_texture[64][32] = 0;	doodle_left_transparency_texture[64][33] = 0;	doodle_left_transparency_texture[64][34] = 0;	doodle_left_transparency_texture[64][35] = 0;	doodle_left_transparency_texture[64][36] = 1;	doodle_left_transparency_texture[64][37] = 1;	doodle_left_transparency_texture[64][38] = 1;	doodle_left_transparency_texture[64][39] = 1;	doodle_left_transparency_texture[64][40] = 1;	doodle_left_transparency_texture[64][41] = 1;	doodle_left_transparency_texture[64][42] = 1;	doodle_left_transparency_texture[64][43] = 1;	doodle_left_transparency_texture[64][44] = 0;	doodle_left_transparency_texture[64][45] = 0;	doodle_left_transparency_texture[64][46] = 0;	doodle_left_transparency_texture[64][47] = 0;	doodle_left_transparency_texture[64][48] = 1;	doodle_left_transparency_texture[64][49] = 1;	doodle_left_transparency_texture[64][50] = 1;	doodle_left_transparency_texture[64][51] = 1;	doodle_left_transparency_texture[64][52] = 1;	doodle_left_transparency_texture[64][53] = 1;	doodle_left_transparency_texture[64][54] = 1;	doodle_left_transparency_texture[64][55] = 1;	doodle_left_transparency_texture[64][56] = 0;	doodle_left_transparency_texture[64][57] = 0;	doodle_left_transparency_texture[64][58] = 0;	doodle_left_transparency_texture[64][59] = 0;	doodle_left_transparency_texture[64][60] = 1;	doodle_left_transparency_texture[64][61] = 1;	doodle_left_transparency_texture[64][62] = 1;	doodle_left_transparency_texture[64][63] = 1;	doodle_left_transparency_texture[64][64] = 1;	doodle_left_transparency_texture[64][65] = 1;	doodle_left_transparency_texture[64][66] = 1;	doodle_left_transparency_texture[64][67] = 1;	doodle_left_transparency_texture[64][68] = 0;	doodle_left_transparency_texture[64][69] = 0;	doodle_left_transparency_texture[64][70] = 0;	doodle_left_transparency_texture[64][71] = 0;	doodle_left_transparency_texture[64][72] = 1;	doodle_left_transparency_texture[64][73] = 1;	doodle_left_transparency_texture[64][74] = 1;	doodle_left_transparency_texture[64][75] = 1;	doodle_left_transparency_texture[64][76] = 1;	doodle_left_transparency_texture[64][77] = 1;	doodle_left_transparency_texture[64][78] = 1;	doodle_left_transparency_texture[64][79] = 1;	doodle_left_transparency_texture[65][0] = 1;	doodle_left_transparency_texture[65][1] = 1;	doodle_left_transparency_texture[65][2] = 1;	doodle_left_transparency_texture[65][3] = 1;	doodle_left_transparency_texture[65][4] = 1;	doodle_left_transparency_texture[65][5] = 1;	doodle_left_transparency_texture[65][6] = 1;	doodle_left_transparency_texture[65][7] = 1;	doodle_left_transparency_texture[65][8] = 1;	doodle_left_transparency_texture[65][9] = 1;	doodle_left_transparency_texture[65][10] = 1;	doodle_left_transparency_texture[65][11] = 1;	doodle_left_transparency_texture[65][12] = 1;	doodle_left_transparency_texture[65][13] = 1;	doodle_left_transparency_texture[65][14] = 1;	doodle_left_transparency_texture[65][15] = 1;	doodle_left_transparency_texture[65][16] = 1;	doodle_left_transparency_texture[65][17] = 1;	doodle_left_transparency_texture[65][18] = 1;	doodle_left_transparency_texture[65][19] = 1;	doodle_left_transparency_texture[65][20] = 1;	doodle_left_transparency_texture[65][21] = 1;	doodle_left_transparency_texture[65][22] = 1;	doodle_left_transparency_texture[65][23] = 1;	doodle_left_transparency_texture[65][24] = 1;	doodle_left_transparency_texture[65][25] = 1;	doodle_left_transparency_texture[65][26] = 1;	doodle_left_transparency_texture[65][27] = 1;	doodle_left_transparency_texture[65][28] = 1;	doodle_left_transparency_texture[65][29] = 1;	doodle_left_transparency_texture[65][30] = 1;	doodle_left_transparency_texture[65][31] = 1;	doodle_left_transparency_texture[65][32] = 0;	doodle_left_transparency_texture[65][33] = 0;	doodle_left_transparency_texture[65][34] = 0;	doodle_left_transparency_texture[65][35] = 0;	doodle_left_transparency_texture[65][36] = 1;	doodle_left_transparency_texture[65][37] = 1;	doodle_left_transparency_texture[65][38] = 1;	doodle_left_transparency_texture[65][39] = 1;	doodle_left_transparency_texture[65][40] = 1;	doodle_left_transparency_texture[65][41] = 1;	doodle_left_transparency_texture[65][42] = 1;	doodle_left_transparency_texture[65][43] = 1;	doodle_left_transparency_texture[65][44] = 0;	doodle_left_transparency_texture[65][45] = 0;	doodle_left_transparency_texture[65][46] = 0;	doodle_left_transparency_texture[65][47] = 0;	doodle_left_transparency_texture[65][48] = 1;	doodle_left_transparency_texture[65][49] = 1;	doodle_left_transparency_texture[65][50] = 1;	doodle_left_transparency_texture[65][51] = 1;	doodle_left_transparency_texture[65][52] = 1;	doodle_left_transparency_texture[65][53] = 1;	doodle_left_transparency_texture[65][54] = 1;	doodle_left_transparency_texture[65][55] = 1;	doodle_left_transparency_texture[65][56] = 0;	doodle_left_transparency_texture[65][57] = 0;	doodle_left_transparency_texture[65][58] = 0;	doodle_left_transparency_texture[65][59] = 0;	doodle_left_transparency_texture[65][60] = 1;	doodle_left_transparency_texture[65][61] = 1;	doodle_left_transparency_texture[65][62] = 1;	doodle_left_transparency_texture[65][63] = 1;	doodle_left_transparency_texture[65][64] = 1;	doodle_left_transparency_texture[65][65] = 1;	doodle_left_transparency_texture[65][66] = 1;	doodle_left_transparency_texture[65][67] = 1;	doodle_left_transparency_texture[65][68] = 0;	doodle_left_transparency_texture[65][69] = 0;	doodle_left_transparency_texture[65][70] = 0;	doodle_left_transparency_texture[65][71] = 0;	doodle_left_transparency_texture[65][72] = 1;	doodle_left_transparency_texture[65][73] = 1;	doodle_left_transparency_texture[65][74] = 1;	doodle_left_transparency_texture[65][75] = 1;	doodle_left_transparency_texture[65][76] = 1;	doodle_left_transparency_texture[65][77] = 1;	doodle_left_transparency_texture[65][78] = 1;	doodle_left_transparency_texture[65][79] = 1;	doodle_left_transparency_texture[66][0] = 1;	doodle_left_transparency_texture[66][1] = 1;	doodle_left_transparency_texture[66][2] = 1;	doodle_left_transparency_texture[66][3] = 1;	doodle_left_transparency_texture[66][4] = 1;	doodle_left_transparency_texture[66][5] = 1;	doodle_left_transparency_texture[66][6] = 1;	doodle_left_transparency_texture[66][7] = 1;	doodle_left_transparency_texture[66][8] = 1;	doodle_left_transparency_texture[66][9] = 1;	doodle_left_transparency_texture[66][10] = 1;	doodle_left_transparency_texture[66][11] = 1;	doodle_left_transparency_texture[66][12] = 1;	doodle_left_transparency_texture[66][13] = 1;	doodle_left_transparency_texture[66][14] = 1;	doodle_left_transparency_texture[66][15] = 1;	doodle_left_transparency_texture[66][16] = 1;	doodle_left_transparency_texture[66][17] = 1;	doodle_left_transparency_texture[66][18] = 1;	doodle_left_transparency_texture[66][19] = 1;	doodle_left_transparency_texture[66][20] = 1;	doodle_left_transparency_texture[66][21] = 1;	doodle_left_transparency_texture[66][22] = 1;	doodle_left_transparency_texture[66][23] = 1;	doodle_left_transparency_texture[66][24] = 1;	doodle_left_transparency_texture[66][25] = 1;	doodle_left_transparency_texture[66][26] = 1;	doodle_left_transparency_texture[66][27] = 1;	doodle_left_transparency_texture[66][28] = 1;	doodle_left_transparency_texture[66][29] = 1;	doodle_left_transparency_texture[66][30] = 1;	doodle_left_transparency_texture[66][31] = 1;	doodle_left_transparency_texture[66][32] = 0;	doodle_left_transparency_texture[66][33] = 0;	doodle_left_transparency_texture[66][34] = 0;	doodle_left_transparency_texture[66][35] = 0;	doodle_left_transparency_texture[66][36] = 1;	doodle_left_transparency_texture[66][37] = 1;	doodle_left_transparency_texture[66][38] = 1;	doodle_left_transparency_texture[66][39] = 1;	doodle_left_transparency_texture[66][40] = 1;	doodle_left_transparency_texture[66][41] = 1;	doodle_left_transparency_texture[66][42] = 1;	doodle_left_transparency_texture[66][43] = 1;	doodle_left_transparency_texture[66][44] = 0;	doodle_left_transparency_texture[66][45] = 0;	doodle_left_transparency_texture[66][46] = 0;	doodle_left_transparency_texture[66][47] = 0;	doodle_left_transparency_texture[66][48] = 1;	doodle_left_transparency_texture[66][49] = 1;	doodle_left_transparency_texture[66][50] = 1;	doodle_left_transparency_texture[66][51] = 1;	doodle_left_transparency_texture[66][52] = 1;	doodle_left_transparency_texture[66][53] = 1;	doodle_left_transparency_texture[66][54] = 1;	doodle_left_transparency_texture[66][55] = 1;	doodle_left_transparency_texture[66][56] = 0;	doodle_left_transparency_texture[66][57] = 0;	doodle_left_transparency_texture[66][58] = 0;	doodle_left_transparency_texture[66][59] = 0;	doodle_left_transparency_texture[66][60] = 1;	doodle_left_transparency_texture[66][61] = 1;	doodle_left_transparency_texture[66][62] = 1;	doodle_left_transparency_texture[66][63] = 1;	doodle_left_transparency_texture[66][64] = 1;	doodle_left_transparency_texture[66][65] = 1;	doodle_left_transparency_texture[66][66] = 1;	doodle_left_transparency_texture[66][67] = 1;	doodle_left_transparency_texture[66][68] = 0;	doodle_left_transparency_texture[66][69] = 0;	doodle_left_transparency_texture[66][70] = 0;	doodle_left_transparency_texture[66][71] = 0;	doodle_left_transparency_texture[66][72] = 1;	doodle_left_transparency_texture[66][73] = 1;	doodle_left_transparency_texture[66][74] = 1;	doodle_left_transparency_texture[66][75] = 1;	doodle_left_transparency_texture[66][76] = 1;	doodle_left_transparency_texture[66][77] = 1;	doodle_left_transparency_texture[66][78] = 1;	doodle_left_transparency_texture[66][79] = 1;	doodle_left_transparency_texture[67][0] = 1;	doodle_left_transparency_texture[67][1] = 1;	doodle_left_transparency_texture[67][2] = 1;	doodle_left_transparency_texture[67][3] = 1;	doodle_left_transparency_texture[67][4] = 1;	doodle_left_transparency_texture[67][5] = 1;	doodle_left_transparency_texture[67][6] = 1;	doodle_left_transparency_texture[67][7] = 1;	doodle_left_transparency_texture[67][8] = 1;	doodle_left_transparency_texture[67][9] = 1;	doodle_left_transparency_texture[67][10] = 1;	doodle_left_transparency_texture[67][11] = 1;	doodle_left_transparency_texture[67][12] = 1;	doodle_left_transparency_texture[67][13] = 1;	doodle_left_transparency_texture[67][14] = 1;	doodle_left_transparency_texture[67][15] = 1;	doodle_left_transparency_texture[67][16] = 1;	doodle_left_transparency_texture[67][17] = 1;	doodle_left_transparency_texture[67][18] = 1;	doodle_left_transparency_texture[67][19] = 1;	doodle_left_transparency_texture[67][20] = 1;	doodle_left_transparency_texture[67][21] = 1;	doodle_left_transparency_texture[67][22] = 1;	doodle_left_transparency_texture[67][23] = 1;	doodle_left_transparency_texture[67][24] = 1;	doodle_left_transparency_texture[67][25] = 1;	doodle_left_transparency_texture[67][26] = 1;	doodle_left_transparency_texture[67][27] = 1;	doodle_left_transparency_texture[67][28] = 1;	doodle_left_transparency_texture[67][29] = 1;	doodle_left_transparency_texture[67][30] = 1;	doodle_left_transparency_texture[67][31] = 1;	doodle_left_transparency_texture[67][32] = 0;	doodle_left_transparency_texture[67][33] = 0;	doodle_left_transparency_texture[67][34] = 0;	doodle_left_transparency_texture[67][35] = 0;	doodle_left_transparency_texture[67][36] = 1;	doodle_left_transparency_texture[67][37] = 1;	doodle_left_transparency_texture[67][38] = 1;	doodle_left_transparency_texture[67][39] = 1;	doodle_left_transparency_texture[67][40] = 1;	doodle_left_transparency_texture[67][41] = 1;	doodle_left_transparency_texture[67][42] = 1;	doodle_left_transparency_texture[67][43] = 1;	doodle_left_transparency_texture[67][44] = 0;	doodle_left_transparency_texture[67][45] = 0;	doodle_left_transparency_texture[67][46] = 0;	doodle_left_transparency_texture[67][47] = 0;	doodle_left_transparency_texture[67][48] = 1;	doodle_left_transparency_texture[67][49] = 1;	doodle_left_transparency_texture[67][50] = 1;	doodle_left_transparency_texture[67][51] = 1;	doodle_left_transparency_texture[67][52] = 1;	doodle_left_transparency_texture[67][53] = 1;	doodle_left_transparency_texture[67][54] = 1;	doodle_left_transparency_texture[67][55] = 1;	doodle_left_transparency_texture[67][56] = 0;	doodle_left_transparency_texture[67][57] = 0;	doodle_left_transparency_texture[67][58] = 0;	doodle_left_transparency_texture[67][59] = 0;	doodle_left_transparency_texture[67][60] = 1;	doodle_left_transparency_texture[67][61] = 1;	doodle_left_transparency_texture[67][62] = 1;	doodle_left_transparency_texture[67][63] = 1;	doodle_left_transparency_texture[67][64] = 1;	doodle_left_transparency_texture[67][65] = 1;	doodle_left_transparency_texture[67][66] = 1;	doodle_left_transparency_texture[67][67] = 1;	doodle_left_transparency_texture[67][68] = 0;	doodle_left_transparency_texture[67][69] = 0;	doodle_left_transparency_texture[67][70] = 0;	doodle_left_transparency_texture[67][71] = 0;	doodle_left_transparency_texture[67][72] = 1;	doodle_left_transparency_texture[67][73] = 1;	doodle_left_transparency_texture[67][74] = 1;	doodle_left_transparency_texture[67][75] = 1;	doodle_left_transparency_texture[67][76] = 1;	doodle_left_transparency_texture[67][77] = 1;	doodle_left_transparency_texture[67][78] = 1;	doodle_left_transparency_texture[67][79] = 1;	doodle_left_transparency_texture[68][0] = 1;	doodle_left_transparency_texture[68][1] = 1;	doodle_left_transparency_texture[68][2] = 1;	doodle_left_transparency_texture[68][3] = 1;	doodle_left_transparency_texture[68][4] = 1;	doodle_left_transparency_texture[68][5] = 1;	doodle_left_transparency_texture[68][6] = 1;	doodle_left_transparency_texture[68][7] = 1;	doodle_left_transparency_texture[68][8] = 1;	doodle_left_transparency_texture[68][9] = 1;	doodle_left_transparency_texture[68][10] = 1;	doodle_left_transparency_texture[68][11] = 1;	doodle_left_transparency_texture[68][12] = 1;	doodle_left_transparency_texture[68][13] = 1;	doodle_left_transparency_texture[68][14] = 1;	doodle_left_transparency_texture[68][15] = 1;	doodle_left_transparency_texture[68][16] = 1;	doodle_left_transparency_texture[68][17] = 1;	doodle_left_transparency_texture[68][18] = 1;	doodle_left_transparency_texture[68][19] = 1;	doodle_left_transparency_texture[68][20] = 1;	doodle_left_transparency_texture[68][21] = 1;	doodle_left_transparency_texture[68][22] = 1;	doodle_left_transparency_texture[68][23] = 1;	doodle_left_transparency_texture[68][24] = 1;	doodle_left_transparency_texture[68][25] = 1;	doodle_left_transparency_texture[68][26] = 1;	doodle_left_transparency_texture[68][27] = 1;	doodle_left_transparency_texture[68][28] = 0;	doodle_left_transparency_texture[68][29] = 0;	doodle_left_transparency_texture[68][30] = 0;	doodle_left_transparency_texture[68][31] = 0;	doodle_left_transparency_texture[68][32] = 0;	doodle_left_transparency_texture[68][33] = 0;	doodle_left_transparency_texture[68][34] = 0;	doodle_left_transparency_texture[68][35] = 0;	doodle_left_transparency_texture[68][36] = 1;	doodle_left_transparency_texture[68][37] = 1;	doodle_left_transparency_texture[68][38] = 1;	doodle_left_transparency_texture[68][39] = 1;	doodle_left_transparency_texture[68][40] = 0;	doodle_left_transparency_texture[68][41] = 0;	doodle_left_transparency_texture[68][42] = 0;	doodle_left_transparency_texture[68][43] = 0;	doodle_left_transparency_texture[68][44] = 0;	doodle_left_transparency_texture[68][45] = 0;	doodle_left_transparency_texture[68][46] = 0;	doodle_left_transparency_texture[68][47] = 0;	doodle_left_transparency_texture[68][48] = 1;	doodle_left_transparency_texture[68][49] = 1;	doodle_left_transparency_texture[68][50] = 1;	doodle_left_transparency_texture[68][51] = 1;	doodle_left_transparency_texture[68][52] = 0;	doodle_left_transparency_texture[68][53] = 0;	doodle_left_transparency_texture[68][54] = 0;	doodle_left_transparency_texture[68][55] = 0;	doodle_left_transparency_texture[68][56] = 0;	doodle_left_transparency_texture[68][57] = 0;	doodle_left_transparency_texture[68][58] = 0;	doodle_left_transparency_texture[68][59] = 0;	doodle_left_transparency_texture[68][60] = 1;	doodle_left_transparency_texture[68][61] = 1;	doodle_left_transparency_texture[68][62] = 1;	doodle_left_transparency_texture[68][63] = 1;	doodle_left_transparency_texture[68][64] = 0;	doodle_left_transparency_texture[68][65] = 0;	doodle_left_transparency_texture[68][66] = 0;	doodle_left_transparency_texture[68][67] = 0;	doodle_left_transparency_texture[68][68] = 0;	doodle_left_transparency_texture[68][69] = 0;	doodle_left_transparency_texture[68][70] = 0;	doodle_left_transparency_texture[68][71] = 0;	doodle_left_transparency_texture[68][72] = 1;	doodle_left_transparency_texture[68][73] = 1;	doodle_left_transparency_texture[68][74] = 1;	doodle_left_transparency_texture[68][75] = 1;	doodle_left_transparency_texture[68][76] = 1;	doodle_left_transparency_texture[68][77] = 1;	doodle_left_transparency_texture[68][78] = 1;	doodle_left_transparency_texture[68][79] = 1;	doodle_left_transparency_texture[69][0] = 1;	doodle_left_transparency_texture[69][1] = 1;	doodle_left_transparency_texture[69][2] = 1;	doodle_left_transparency_texture[69][3] = 1;	doodle_left_transparency_texture[69][4] = 1;	doodle_left_transparency_texture[69][5] = 1;	doodle_left_transparency_texture[69][6] = 1;	doodle_left_transparency_texture[69][7] = 1;	doodle_left_transparency_texture[69][8] = 1;	doodle_left_transparency_texture[69][9] = 1;	doodle_left_transparency_texture[69][10] = 1;	doodle_left_transparency_texture[69][11] = 1;	doodle_left_transparency_texture[69][12] = 1;	doodle_left_transparency_texture[69][13] = 1;	doodle_left_transparency_texture[69][14] = 1;	doodle_left_transparency_texture[69][15] = 1;	doodle_left_transparency_texture[69][16] = 1;	doodle_left_transparency_texture[69][17] = 1;	doodle_left_transparency_texture[69][18] = 1;	doodle_left_transparency_texture[69][19] = 1;	doodle_left_transparency_texture[69][20] = 1;	doodle_left_transparency_texture[69][21] = 1;	doodle_left_transparency_texture[69][22] = 1;	doodle_left_transparency_texture[69][23] = 1;	doodle_left_transparency_texture[69][24] = 1;	doodle_left_transparency_texture[69][25] = 1;	doodle_left_transparency_texture[69][26] = 1;	doodle_left_transparency_texture[69][27] = 1;	doodle_left_transparency_texture[69][28] = 0;	doodle_left_transparency_texture[69][29] = 0;	doodle_left_transparency_texture[69][30] = 0;	doodle_left_transparency_texture[69][31] = 0;	doodle_left_transparency_texture[69][32] = 0;	doodle_left_transparency_texture[69][33] = 0;	doodle_left_transparency_texture[69][34] = 0;	doodle_left_transparency_texture[69][35] = 0;	doodle_left_transparency_texture[69][36] = 1;	doodle_left_transparency_texture[69][37] = 1;	doodle_left_transparency_texture[69][38] = 1;	doodle_left_transparency_texture[69][39] = 1;	doodle_left_transparency_texture[69][40] = 0;	doodle_left_transparency_texture[69][41] = 0;	doodle_left_transparency_texture[69][42] = 0;	doodle_left_transparency_texture[69][43] = 0;	doodle_left_transparency_texture[69][44] = 0;	doodle_left_transparency_texture[69][45] = 0;	doodle_left_transparency_texture[69][46] = 0;	doodle_left_transparency_texture[69][47] = 0;	doodle_left_transparency_texture[69][48] = 1;	doodle_left_transparency_texture[69][49] = 1;	doodle_left_transparency_texture[69][50] = 1;	doodle_left_transparency_texture[69][51] = 1;	doodle_left_transparency_texture[69][52] = 0;	doodle_left_transparency_texture[69][53] = 0;	doodle_left_transparency_texture[69][54] = 0;	doodle_left_transparency_texture[69][55] = 0;	doodle_left_transparency_texture[69][56] = 0;	doodle_left_transparency_texture[69][57] = 0;	doodle_left_transparency_texture[69][58] = 0;	doodle_left_transparency_texture[69][59] = 0;	doodle_left_transparency_texture[69][60] = 1;	doodle_left_transparency_texture[69][61] = 1;	doodle_left_transparency_texture[69][62] = 1;	doodle_left_transparency_texture[69][63] = 1;	doodle_left_transparency_texture[69][64] = 0;	doodle_left_transparency_texture[69][65] = 0;	doodle_left_transparency_texture[69][66] = 0;	doodle_left_transparency_texture[69][67] = 0;	doodle_left_transparency_texture[69][68] = 0;	doodle_left_transparency_texture[69][69] = 0;	doodle_left_transparency_texture[69][70] = 0;	doodle_left_transparency_texture[69][71] = 0;	doodle_left_transparency_texture[69][72] = 1;	doodle_left_transparency_texture[69][73] = 1;	doodle_left_transparency_texture[69][74] = 1;	doodle_left_transparency_texture[69][75] = 1;	doodle_left_transparency_texture[69][76] = 1;	doodle_left_transparency_texture[69][77] = 1;	doodle_left_transparency_texture[69][78] = 1;	doodle_left_transparency_texture[69][79] = 1;	doodle_left_transparency_texture[70][0] = 1;	doodle_left_transparency_texture[70][1] = 1;	doodle_left_transparency_texture[70][2] = 1;	doodle_left_transparency_texture[70][3] = 1;	doodle_left_transparency_texture[70][4] = 1;	doodle_left_transparency_texture[70][5] = 1;	doodle_left_transparency_texture[70][6] = 1;	doodle_left_transparency_texture[70][7] = 1;	doodle_left_transparency_texture[70][8] = 1;	doodle_left_transparency_texture[70][9] = 1;	doodle_left_transparency_texture[70][10] = 1;	doodle_left_transparency_texture[70][11] = 1;	doodle_left_transparency_texture[70][12] = 1;	doodle_left_transparency_texture[70][13] = 1;	doodle_left_transparency_texture[70][14] = 1;	doodle_left_transparency_texture[70][15] = 1;	doodle_left_transparency_texture[70][16] = 1;	doodle_left_transparency_texture[70][17] = 1;	doodle_left_transparency_texture[70][18] = 1;	doodle_left_transparency_texture[70][19] = 1;	doodle_left_transparency_texture[70][20] = 1;	doodle_left_transparency_texture[70][21] = 1;	doodle_left_transparency_texture[70][22] = 1;	doodle_left_transparency_texture[70][23] = 1;	doodle_left_transparency_texture[70][24] = 1;	doodle_left_transparency_texture[70][25] = 1;	doodle_left_transparency_texture[70][26] = 1;	doodle_left_transparency_texture[70][27] = 1;	doodle_left_transparency_texture[70][28] = 0;	doodle_left_transparency_texture[70][29] = 0;	doodle_left_transparency_texture[70][30] = 0;	doodle_left_transparency_texture[70][31] = 0;	doodle_left_transparency_texture[70][32] = 0;	doodle_left_transparency_texture[70][33] = 0;	doodle_left_transparency_texture[70][34] = 0;	doodle_left_transparency_texture[70][35] = 0;	doodle_left_transparency_texture[70][36] = 1;	doodle_left_transparency_texture[70][37] = 1;	doodle_left_transparency_texture[70][38] = 1;	doodle_left_transparency_texture[70][39] = 1;	doodle_left_transparency_texture[70][40] = 0;	doodle_left_transparency_texture[70][41] = 0;	doodle_left_transparency_texture[70][42] = 0;	doodle_left_transparency_texture[70][43] = 0;	doodle_left_transparency_texture[70][44] = 0;	doodle_left_transparency_texture[70][45] = 0;	doodle_left_transparency_texture[70][46] = 0;	doodle_left_transparency_texture[70][47] = 0;	doodle_left_transparency_texture[70][48] = 1;	doodle_left_transparency_texture[70][49] = 1;	doodle_left_transparency_texture[70][50] = 1;	doodle_left_transparency_texture[70][51] = 1;	doodle_left_transparency_texture[70][52] = 0;	doodle_left_transparency_texture[70][53] = 0;	doodle_left_transparency_texture[70][54] = 0;	doodle_left_transparency_texture[70][55] = 0;	doodle_left_transparency_texture[70][56] = 0;	doodle_left_transparency_texture[70][57] = 0;	doodle_left_transparency_texture[70][58] = 0;	doodle_left_transparency_texture[70][59] = 0;	doodle_left_transparency_texture[70][60] = 1;	doodle_left_transparency_texture[70][61] = 1;	doodle_left_transparency_texture[70][62] = 1;	doodle_left_transparency_texture[70][63] = 1;	doodle_left_transparency_texture[70][64] = 0;	doodle_left_transparency_texture[70][65] = 0;	doodle_left_transparency_texture[70][66] = 0;	doodle_left_transparency_texture[70][67] = 0;	doodle_left_transparency_texture[70][68] = 0;	doodle_left_transparency_texture[70][69] = 0;	doodle_left_transparency_texture[70][70] = 0;	doodle_left_transparency_texture[70][71] = 0;	doodle_left_transparency_texture[70][72] = 1;	doodle_left_transparency_texture[70][73] = 1;	doodle_left_transparency_texture[70][74] = 1;	doodle_left_transparency_texture[70][75] = 1;	doodle_left_transparency_texture[70][76] = 1;	doodle_left_transparency_texture[70][77] = 1;	doodle_left_transparency_texture[70][78] = 1;	doodle_left_transparency_texture[70][79] = 1;	doodle_left_transparency_texture[71][0] = 1;	doodle_left_transparency_texture[71][1] = 1;	doodle_left_transparency_texture[71][2] = 1;	doodle_left_transparency_texture[71][3] = 1;	doodle_left_transparency_texture[71][4] = 1;	doodle_left_transparency_texture[71][5] = 1;	doodle_left_transparency_texture[71][6] = 1;	doodle_left_transparency_texture[71][7] = 1;	doodle_left_transparency_texture[71][8] = 1;	doodle_left_transparency_texture[71][9] = 1;	doodle_left_transparency_texture[71][10] = 1;	doodle_left_transparency_texture[71][11] = 1;	doodle_left_transparency_texture[71][12] = 1;	doodle_left_transparency_texture[71][13] = 1;	doodle_left_transparency_texture[71][14] = 1;	doodle_left_transparency_texture[71][15] = 1;	doodle_left_transparency_texture[71][16] = 1;	doodle_left_transparency_texture[71][17] = 1;	doodle_left_transparency_texture[71][18] = 1;	doodle_left_transparency_texture[71][19] = 1;	doodle_left_transparency_texture[71][20] = 1;	doodle_left_transparency_texture[71][21] = 1;	doodle_left_transparency_texture[71][22] = 1;	doodle_left_transparency_texture[71][23] = 1;	doodle_left_transparency_texture[71][24] = 1;	doodle_left_transparency_texture[71][25] = 1;	doodle_left_transparency_texture[71][26] = 1;	doodle_left_transparency_texture[71][27] = 1;	doodle_left_transparency_texture[71][28] = 0;	doodle_left_transparency_texture[71][29] = 0;	doodle_left_transparency_texture[71][30] = 0;	doodle_left_transparency_texture[71][31] = 0;	doodle_left_transparency_texture[71][32] = 0;	doodle_left_transparency_texture[71][33] = 0;	doodle_left_transparency_texture[71][34] = 0;	doodle_left_transparency_texture[71][35] = 0;	doodle_left_transparency_texture[71][36] = 1;	doodle_left_transparency_texture[71][37] = 1;	doodle_left_transparency_texture[71][38] = 1;	doodle_left_transparency_texture[71][39] = 1;	doodle_left_transparency_texture[71][40] = 0;	doodle_left_transparency_texture[71][41] = 0;	doodle_left_transparency_texture[71][42] = 0;	doodle_left_transparency_texture[71][43] = 0;	doodle_left_transparency_texture[71][44] = 0;	doodle_left_transparency_texture[71][45] = 0;	doodle_left_transparency_texture[71][46] = 0;	doodle_left_transparency_texture[71][47] = 0;	doodle_left_transparency_texture[71][48] = 1;	doodle_left_transparency_texture[71][49] = 1;	doodle_left_transparency_texture[71][50] = 1;	doodle_left_transparency_texture[71][51] = 1;	doodle_left_transparency_texture[71][52] = 0;	doodle_left_transparency_texture[71][53] = 0;	doodle_left_transparency_texture[71][54] = 0;	doodle_left_transparency_texture[71][55] = 0;	doodle_left_transparency_texture[71][56] = 0;	doodle_left_transparency_texture[71][57] = 0;	doodle_left_transparency_texture[71][58] = 0;	doodle_left_transparency_texture[71][59] = 0;	doodle_left_transparency_texture[71][60] = 1;	doodle_left_transparency_texture[71][61] = 1;	doodle_left_transparency_texture[71][62] = 1;	doodle_left_transparency_texture[71][63] = 1;	doodle_left_transparency_texture[71][64] = 0;	doodle_left_transparency_texture[71][65] = 0;	doodle_left_transparency_texture[71][66] = 0;	doodle_left_transparency_texture[71][67] = 0;	doodle_left_transparency_texture[71][68] = 0;	doodle_left_transparency_texture[71][69] = 0;	doodle_left_transparency_texture[71][70] = 0;	doodle_left_transparency_texture[71][71] = 0;	doodle_left_transparency_texture[71][72] = 1;	doodle_left_transparency_texture[71][73] = 1;	doodle_left_transparency_texture[71][74] = 1;	doodle_left_transparency_texture[71][75] = 1;	doodle_left_transparency_texture[71][76] = 1;	doodle_left_transparency_texture[71][77] = 1;	doodle_left_transparency_texture[71][78] = 1;	doodle_left_transparency_texture[71][79] = 1;	doodle_left_transparency_texture[72][0] = 1;	doodle_left_transparency_texture[72][1] = 1;	doodle_left_transparency_texture[72][2] = 1;	doodle_left_transparency_texture[72][3] = 1;	doodle_left_transparency_texture[72][4] = 1;	doodle_left_transparency_texture[72][5] = 1;	doodle_left_transparency_texture[72][6] = 1;	doodle_left_transparency_texture[72][7] = 1;	doodle_left_transparency_texture[72][8] = 1;	doodle_left_transparency_texture[72][9] = 1;	doodle_left_transparency_texture[72][10] = 1;	doodle_left_transparency_texture[72][11] = 1;	doodle_left_transparency_texture[72][12] = 1;	doodle_left_transparency_texture[72][13] = 1;	doodle_left_transparency_texture[72][14] = 1;	doodle_left_transparency_texture[72][15] = 1;	doodle_left_transparency_texture[72][16] = 1;	doodle_left_transparency_texture[72][17] = 1;	doodle_left_transparency_texture[72][18] = 1;	doodle_left_transparency_texture[72][19] = 1;	doodle_left_transparency_texture[72][20] = 1;	doodle_left_transparency_texture[72][21] = 1;	doodle_left_transparency_texture[72][22] = 1;	doodle_left_transparency_texture[72][23] = 1;	doodle_left_transparency_texture[72][24] = 1;	doodle_left_transparency_texture[72][25] = 1;	doodle_left_transparency_texture[72][26] = 1;	doodle_left_transparency_texture[72][27] = 1;	doodle_left_transparency_texture[72][28] = 1;	doodle_left_transparency_texture[72][29] = 1;	doodle_left_transparency_texture[72][30] = 1;	doodle_left_transparency_texture[72][31] = 1;	doodle_left_transparency_texture[72][32] = 1;	doodle_left_transparency_texture[72][33] = 1;	doodle_left_transparency_texture[72][34] = 1;	doodle_left_transparency_texture[72][35] = 1;	doodle_left_transparency_texture[72][36] = 1;	doodle_left_transparency_texture[72][37] = 1;	doodle_left_transparency_texture[72][38] = 1;	doodle_left_transparency_texture[72][39] = 1;	doodle_left_transparency_texture[72][40] = 1;	doodle_left_transparency_texture[72][41] = 1;	doodle_left_transparency_texture[72][42] = 1;	doodle_left_transparency_texture[72][43] = 1;	doodle_left_transparency_texture[72][44] = 1;	doodle_left_transparency_texture[72][45] = 1;	doodle_left_transparency_texture[72][46] = 1;	doodle_left_transparency_texture[72][47] = 1;	doodle_left_transparency_texture[72][48] = 1;	doodle_left_transparency_texture[72][49] = 1;	doodle_left_transparency_texture[72][50] = 1;	doodle_left_transparency_texture[72][51] = 1;	doodle_left_transparency_texture[72][52] = 1;	doodle_left_transparency_texture[72][53] = 1;	doodle_left_transparency_texture[72][54] = 1;	doodle_left_transparency_texture[72][55] = 1;	doodle_left_transparency_texture[72][56] = 1;	doodle_left_transparency_texture[72][57] = 1;	doodle_left_transparency_texture[72][58] = 1;	doodle_left_transparency_texture[72][59] = 1;	doodle_left_transparency_texture[72][60] = 1;	doodle_left_transparency_texture[72][61] = 1;	doodle_left_transparency_texture[72][62] = 1;	doodle_left_transparency_texture[72][63] = 1;	doodle_left_transparency_texture[72][64] = 1;	doodle_left_transparency_texture[72][65] = 1;	doodle_left_transparency_texture[72][66] = 1;	doodle_left_transparency_texture[72][67] = 1;	doodle_left_transparency_texture[72][68] = 1;	doodle_left_transparency_texture[72][69] = 1;	doodle_left_transparency_texture[72][70] = 1;	doodle_left_transparency_texture[72][71] = 1;	doodle_left_transparency_texture[72][72] = 1;	doodle_left_transparency_texture[72][73] = 1;	doodle_left_transparency_texture[72][74] = 1;	doodle_left_transparency_texture[72][75] = 1;	doodle_left_transparency_texture[72][76] = 1;	doodle_left_transparency_texture[72][77] = 1;	doodle_left_transparency_texture[72][78] = 1;	doodle_left_transparency_texture[72][79] = 1;	doodle_left_transparency_texture[73][0] = 1;	doodle_left_transparency_texture[73][1] = 1;	doodle_left_transparency_texture[73][2] = 1;	doodle_left_transparency_texture[73][3] = 1;	doodle_left_transparency_texture[73][4] = 1;	doodle_left_transparency_texture[73][5] = 1;	doodle_left_transparency_texture[73][6] = 1;	doodle_left_transparency_texture[73][7] = 1;	doodle_left_transparency_texture[73][8] = 1;	doodle_left_transparency_texture[73][9] = 1;	doodle_left_transparency_texture[73][10] = 1;	doodle_left_transparency_texture[73][11] = 1;	doodle_left_transparency_texture[73][12] = 1;	doodle_left_transparency_texture[73][13] = 1;	doodle_left_transparency_texture[73][14] = 1;	doodle_left_transparency_texture[73][15] = 1;	doodle_left_transparency_texture[73][16] = 1;	doodle_left_transparency_texture[73][17] = 1;	doodle_left_transparency_texture[73][18] = 1;	doodle_left_transparency_texture[73][19] = 1;	doodle_left_transparency_texture[73][20] = 1;	doodle_left_transparency_texture[73][21] = 1;	doodle_left_transparency_texture[73][22] = 1;	doodle_left_transparency_texture[73][23] = 1;	doodle_left_transparency_texture[73][24] = 1;	doodle_left_transparency_texture[73][25] = 1;	doodle_left_transparency_texture[73][26] = 1;	doodle_left_transparency_texture[73][27] = 1;	doodle_left_transparency_texture[73][28] = 1;	doodle_left_transparency_texture[73][29] = 1;	doodle_left_transparency_texture[73][30] = 1;	doodle_left_transparency_texture[73][31] = 1;	doodle_left_transparency_texture[73][32] = 1;	doodle_left_transparency_texture[73][33] = 1;	doodle_left_transparency_texture[73][34] = 1;	doodle_left_transparency_texture[73][35] = 1;	doodle_left_transparency_texture[73][36] = 1;	doodle_left_transparency_texture[73][37] = 1;	doodle_left_transparency_texture[73][38] = 1;	doodle_left_transparency_texture[73][39] = 1;	doodle_left_transparency_texture[73][40] = 1;	doodle_left_transparency_texture[73][41] = 1;	doodle_left_transparency_texture[73][42] = 1;	doodle_left_transparency_texture[73][43] = 1;	doodle_left_transparency_texture[73][44] = 1;	doodle_left_transparency_texture[73][45] = 1;	doodle_left_transparency_texture[73][46] = 1;	doodle_left_transparency_texture[73][47] = 1;	doodle_left_transparency_texture[73][48] = 1;	doodle_left_transparency_texture[73][49] = 1;	doodle_left_transparency_texture[73][50] = 1;	doodle_left_transparency_texture[73][51] = 1;	doodle_left_transparency_texture[73][52] = 1;	doodle_left_transparency_texture[73][53] = 1;	doodle_left_transparency_texture[73][54] = 1;	doodle_left_transparency_texture[73][55] = 1;	doodle_left_transparency_texture[73][56] = 1;	doodle_left_transparency_texture[73][57] = 1;	doodle_left_transparency_texture[73][58] = 1;	doodle_left_transparency_texture[73][59] = 1;	doodle_left_transparency_texture[73][60] = 1;	doodle_left_transparency_texture[73][61] = 1;	doodle_left_transparency_texture[73][62] = 1;	doodle_left_transparency_texture[73][63] = 1;	doodle_left_transparency_texture[73][64] = 1;	doodle_left_transparency_texture[73][65] = 1;	doodle_left_transparency_texture[73][66] = 1;	doodle_left_transparency_texture[73][67] = 1;	doodle_left_transparency_texture[73][68] = 1;	doodle_left_transparency_texture[73][69] = 1;	doodle_left_transparency_texture[73][70] = 1;	doodle_left_transparency_texture[73][71] = 1;	doodle_left_transparency_texture[73][72] = 1;	doodle_left_transparency_texture[73][73] = 1;	doodle_left_transparency_texture[73][74] = 1;	doodle_left_transparency_texture[73][75] = 1;	doodle_left_transparency_texture[73][76] = 1;	doodle_left_transparency_texture[73][77] = 1;	doodle_left_transparency_texture[73][78] = 1;	doodle_left_transparency_texture[73][79] = 1;	doodle_left_transparency_texture[74][0] = 1;	doodle_left_transparency_texture[74][1] = 1;	doodle_left_transparency_texture[74][2] = 1;	doodle_left_transparency_texture[74][3] = 1;	doodle_left_transparency_texture[74][4] = 1;	doodle_left_transparency_texture[74][5] = 1;	doodle_left_transparency_texture[74][6] = 1;	doodle_left_transparency_texture[74][7] = 1;	doodle_left_transparency_texture[74][8] = 1;	doodle_left_transparency_texture[74][9] = 1;	doodle_left_transparency_texture[74][10] = 1;	doodle_left_transparency_texture[74][11] = 1;	doodle_left_transparency_texture[74][12] = 1;	doodle_left_transparency_texture[74][13] = 1;	doodle_left_transparency_texture[74][14] = 1;	doodle_left_transparency_texture[74][15] = 1;	doodle_left_transparency_texture[74][16] = 1;	doodle_left_transparency_texture[74][17] = 1;	doodle_left_transparency_texture[74][18] = 1;	doodle_left_transparency_texture[74][19] = 1;	doodle_left_transparency_texture[74][20] = 1;	doodle_left_transparency_texture[74][21] = 1;	doodle_left_transparency_texture[74][22] = 1;	doodle_left_transparency_texture[74][23] = 1;	doodle_left_transparency_texture[74][24] = 1;	doodle_left_transparency_texture[74][25] = 1;	doodle_left_transparency_texture[74][26] = 1;	doodle_left_transparency_texture[74][27] = 1;	doodle_left_transparency_texture[74][28] = 1;	doodle_left_transparency_texture[74][29] = 1;	doodle_left_transparency_texture[74][30] = 1;	doodle_left_transparency_texture[74][31] = 1;	doodle_left_transparency_texture[74][32] = 1;	doodle_left_transparency_texture[74][33] = 1;	doodle_left_transparency_texture[74][34] = 1;	doodle_left_transparency_texture[74][35] = 1;	doodle_left_transparency_texture[74][36] = 1;	doodle_left_transparency_texture[74][37] = 1;	doodle_left_transparency_texture[74][38] = 1;	doodle_left_transparency_texture[74][39] = 1;	doodle_left_transparency_texture[74][40] = 1;	doodle_left_transparency_texture[74][41] = 1;	doodle_left_transparency_texture[74][42] = 1;	doodle_left_transparency_texture[74][43] = 1;	doodle_left_transparency_texture[74][44] = 1;	doodle_left_transparency_texture[74][45] = 1;	doodle_left_transparency_texture[74][46] = 1;	doodle_left_transparency_texture[74][47] = 1;	doodle_left_transparency_texture[74][48] = 1;	doodle_left_transparency_texture[74][49] = 1;	doodle_left_transparency_texture[74][50] = 1;	doodle_left_transparency_texture[74][51] = 1;	doodle_left_transparency_texture[74][52] = 1;	doodle_left_transparency_texture[74][53] = 1;	doodle_left_transparency_texture[74][54] = 1;	doodle_left_transparency_texture[74][55] = 1;	doodle_left_transparency_texture[74][56] = 1;	doodle_left_transparency_texture[74][57] = 1;	doodle_left_transparency_texture[74][58] = 1;	doodle_left_transparency_texture[74][59] = 1;	doodle_left_transparency_texture[74][60] = 1;	doodle_left_transparency_texture[74][61] = 1;	doodle_left_transparency_texture[74][62] = 1;	doodle_left_transparency_texture[74][63] = 1;	doodle_left_transparency_texture[74][64] = 1;	doodle_left_transparency_texture[74][65] = 1;	doodle_left_transparency_texture[74][66] = 1;	doodle_left_transparency_texture[74][67] = 1;	doodle_left_transparency_texture[74][68] = 1;	doodle_left_transparency_texture[74][69] = 1;	doodle_left_transparency_texture[74][70] = 1;	doodle_left_transparency_texture[74][71] = 1;	doodle_left_transparency_texture[74][72] = 1;	doodle_left_transparency_texture[74][73] = 1;	doodle_left_transparency_texture[74][74] = 1;	doodle_left_transparency_texture[74][75] = 1;	doodle_left_transparency_texture[74][76] = 1;	doodle_left_transparency_texture[74][77] = 1;	doodle_left_transparency_texture[74][78] = 1;	doodle_left_transparency_texture[74][79] = 1;	doodle_left_transparency_texture[75][0] = 1;	doodle_left_transparency_texture[75][1] = 1;	doodle_left_transparency_texture[75][2] = 1;	doodle_left_transparency_texture[75][3] = 1;	doodle_left_transparency_texture[75][4] = 1;	doodle_left_transparency_texture[75][5] = 1;	doodle_left_transparency_texture[75][6] = 1;	doodle_left_transparency_texture[75][7] = 1;	doodle_left_transparency_texture[75][8] = 1;	doodle_left_transparency_texture[75][9] = 1;	doodle_left_transparency_texture[75][10] = 1;	doodle_left_transparency_texture[75][11] = 1;	doodle_left_transparency_texture[75][12] = 1;	doodle_left_transparency_texture[75][13] = 1;	doodle_left_transparency_texture[75][14] = 1;	doodle_left_transparency_texture[75][15] = 1;	doodle_left_transparency_texture[75][16] = 1;	doodle_left_transparency_texture[75][17] = 1;	doodle_left_transparency_texture[75][18] = 1;	doodle_left_transparency_texture[75][19] = 1;	doodle_left_transparency_texture[75][20] = 1;	doodle_left_transparency_texture[75][21] = 1;	doodle_left_transparency_texture[75][22] = 1;	doodle_left_transparency_texture[75][23] = 1;	doodle_left_transparency_texture[75][24] = 1;	doodle_left_transparency_texture[75][25] = 1;	doodle_left_transparency_texture[75][26] = 1;	doodle_left_transparency_texture[75][27] = 1;	doodle_left_transparency_texture[75][28] = 1;	doodle_left_transparency_texture[75][29] = 1;	doodle_left_transparency_texture[75][30] = 1;	doodle_left_transparency_texture[75][31] = 1;	doodle_left_transparency_texture[75][32] = 1;	doodle_left_transparency_texture[75][33] = 1;	doodle_left_transparency_texture[75][34] = 1;	doodle_left_transparency_texture[75][35] = 1;	doodle_left_transparency_texture[75][36] = 1;	doodle_left_transparency_texture[75][37] = 1;	doodle_left_transparency_texture[75][38] = 1;	doodle_left_transparency_texture[75][39] = 1;	doodle_left_transparency_texture[75][40] = 1;	doodle_left_transparency_texture[75][41] = 1;	doodle_left_transparency_texture[75][42] = 1;	doodle_left_transparency_texture[75][43] = 1;	doodle_left_transparency_texture[75][44] = 1;	doodle_left_transparency_texture[75][45] = 1;	doodle_left_transparency_texture[75][46] = 1;	doodle_left_transparency_texture[75][47] = 1;	doodle_left_transparency_texture[75][48] = 1;	doodle_left_transparency_texture[75][49] = 1;	doodle_left_transparency_texture[75][50] = 1;	doodle_left_transparency_texture[75][51] = 1;	doodle_left_transparency_texture[75][52] = 1;	doodle_left_transparency_texture[75][53] = 1;	doodle_left_transparency_texture[75][54] = 1;	doodle_left_transparency_texture[75][55] = 1;	doodle_left_transparency_texture[75][56] = 1;	doodle_left_transparency_texture[75][57] = 1;	doodle_left_transparency_texture[75][58] = 1;	doodle_left_transparency_texture[75][59] = 1;	doodle_left_transparency_texture[75][60] = 1;	doodle_left_transparency_texture[75][61] = 1;	doodle_left_transparency_texture[75][62] = 1;	doodle_left_transparency_texture[75][63] = 1;	doodle_left_transparency_texture[75][64] = 1;	doodle_left_transparency_texture[75][65] = 1;	doodle_left_transparency_texture[75][66] = 1;	doodle_left_transparency_texture[75][67] = 1;	doodle_left_transparency_texture[75][68] = 1;	doodle_left_transparency_texture[75][69] = 1;	doodle_left_transparency_texture[75][70] = 1;	doodle_left_transparency_texture[75][71] = 1;	doodle_left_transparency_texture[75][72] = 1;	doodle_left_transparency_texture[75][73] = 1;	doodle_left_transparency_texture[75][74] = 1;	doodle_left_transparency_texture[75][75] = 1;	doodle_left_transparency_texture[75][76] = 1;	doodle_left_transparency_texture[75][77] = 1;	doodle_left_transparency_texture[75][78] = 1;	doodle_left_transparency_texture[75][79] = 1;	doodle_left_transparency_texture[76][0] = 1;	doodle_left_transparency_texture[76][1] = 1;	doodle_left_transparency_texture[76][2] = 1;	doodle_left_transparency_texture[76][3] = 1;	doodle_left_transparency_texture[76][4] = 1;	doodle_left_transparency_texture[76][5] = 1;	doodle_left_transparency_texture[76][6] = 1;	doodle_left_transparency_texture[76][7] = 1;	doodle_left_transparency_texture[76][8] = 1;	doodle_left_transparency_texture[76][9] = 1;	doodle_left_transparency_texture[76][10] = 1;	doodle_left_transparency_texture[76][11] = 1;	doodle_left_transparency_texture[76][12] = 1;	doodle_left_transparency_texture[76][13] = 1;	doodle_left_transparency_texture[76][14] = 1;	doodle_left_transparency_texture[76][15] = 1;	doodle_left_transparency_texture[76][16] = 1;	doodle_left_transparency_texture[76][17] = 1;	doodle_left_transparency_texture[76][18] = 1;	doodle_left_transparency_texture[76][19] = 1;	doodle_left_transparency_texture[76][20] = 1;	doodle_left_transparency_texture[76][21] = 1;	doodle_left_transparency_texture[76][22] = 1;	doodle_left_transparency_texture[76][23] = 1;	doodle_left_transparency_texture[76][24] = 1;	doodle_left_transparency_texture[76][25] = 1;	doodle_left_transparency_texture[76][26] = 1;	doodle_left_transparency_texture[76][27] = 1;	doodle_left_transparency_texture[76][28] = 1;	doodle_left_transparency_texture[76][29] = 1;	doodle_left_transparency_texture[76][30] = 1;	doodle_left_transparency_texture[76][31] = 1;	doodle_left_transparency_texture[76][32] = 1;	doodle_left_transparency_texture[76][33] = 1;	doodle_left_transparency_texture[76][34] = 1;	doodle_left_transparency_texture[76][35] = 1;	doodle_left_transparency_texture[76][36] = 1;	doodle_left_transparency_texture[76][37] = 1;	doodle_left_transparency_texture[76][38] = 1;	doodle_left_transparency_texture[76][39] = 1;	doodle_left_transparency_texture[76][40] = 1;	doodle_left_transparency_texture[76][41] = 1;	doodle_left_transparency_texture[76][42] = 1;	doodle_left_transparency_texture[76][43] = 1;	doodle_left_transparency_texture[76][44] = 1;	doodle_left_transparency_texture[76][45] = 1;	doodle_left_transparency_texture[76][46] = 1;	doodle_left_transparency_texture[76][47] = 1;	doodle_left_transparency_texture[76][48] = 1;	doodle_left_transparency_texture[76][49] = 1;	doodle_left_transparency_texture[76][50] = 1;	doodle_left_transparency_texture[76][51] = 1;	doodle_left_transparency_texture[76][52] = 1;	doodle_left_transparency_texture[76][53] = 1;	doodle_left_transparency_texture[76][54] = 1;	doodle_left_transparency_texture[76][55] = 1;	doodle_left_transparency_texture[76][56] = 1;	doodle_left_transparency_texture[76][57] = 1;	doodle_left_transparency_texture[76][58] = 1;	doodle_left_transparency_texture[76][59] = 1;	doodle_left_transparency_texture[76][60] = 1;	doodle_left_transparency_texture[76][61] = 1;	doodle_left_transparency_texture[76][62] = 1;	doodle_left_transparency_texture[76][63] = 1;	doodle_left_transparency_texture[76][64] = 1;	doodle_left_transparency_texture[76][65] = 1;	doodle_left_transparency_texture[76][66] = 1;	doodle_left_transparency_texture[76][67] = 1;	doodle_left_transparency_texture[76][68] = 1;	doodle_left_transparency_texture[76][69] = 1;	doodle_left_transparency_texture[76][70] = 1;	doodle_left_transparency_texture[76][71] = 1;	doodle_left_transparency_texture[76][72] = 1;	doodle_left_transparency_texture[76][73] = 1;	doodle_left_transparency_texture[76][74] = 1;	doodle_left_transparency_texture[76][75] = 1;	doodle_left_transparency_texture[76][76] = 1;	doodle_left_transparency_texture[76][77] = 1;	doodle_left_transparency_texture[76][78] = 1;	doodle_left_transparency_texture[76][79] = 1;	doodle_left_transparency_texture[77][0] = 1;	doodle_left_transparency_texture[77][1] = 1;	doodle_left_transparency_texture[77][2] = 1;	doodle_left_transparency_texture[77][3] = 1;	doodle_left_transparency_texture[77][4] = 1;	doodle_left_transparency_texture[77][5] = 1;	doodle_left_transparency_texture[77][6] = 1;	doodle_left_transparency_texture[77][7] = 1;	doodle_left_transparency_texture[77][8] = 1;	doodle_left_transparency_texture[77][9] = 1;	doodle_left_transparency_texture[77][10] = 1;	doodle_left_transparency_texture[77][11] = 1;	doodle_left_transparency_texture[77][12] = 1;	doodle_left_transparency_texture[77][13] = 1;	doodle_left_transparency_texture[77][14] = 1;	doodle_left_transparency_texture[77][15] = 1;	doodle_left_transparency_texture[77][16] = 1;	doodle_left_transparency_texture[77][17] = 1;	doodle_left_transparency_texture[77][18] = 1;	doodle_left_transparency_texture[77][19] = 1;	doodle_left_transparency_texture[77][20] = 1;	doodle_left_transparency_texture[77][21] = 1;	doodle_left_transparency_texture[77][22] = 1;	doodle_left_transparency_texture[77][23] = 1;	doodle_left_transparency_texture[77][24] = 1;	doodle_left_transparency_texture[77][25] = 1;	doodle_left_transparency_texture[77][26] = 1;	doodle_left_transparency_texture[77][27] = 1;	doodle_left_transparency_texture[77][28] = 1;	doodle_left_transparency_texture[77][29] = 1;	doodle_left_transparency_texture[77][30] = 1;	doodle_left_transparency_texture[77][31] = 1;	doodle_left_transparency_texture[77][32] = 1;	doodle_left_transparency_texture[77][33] = 1;	doodle_left_transparency_texture[77][34] = 1;	doodle_left_transparency_texture[77][35] = 1;	doodle_left_transparency_texture[77][36] = 1;	doodle_left_transparency_texture[77][37] = 1;	doodle_left_transparency_texture[77][38] = 1;	doodle_left_transparency_texture[77][39] = 1;	doodle_left_transparency_texture[77][40] = 1;	doodle_left_transparency_texture[77][41] = 1;	doodle_left_transparency_texture[77][42] = 1;	doodle_left_transparency_texture[77][43] = 1;	doodle_left_transparency_texture[77][44] = 1;	doodle_left_transparency_texture[77][45] = 1;	doodle_left_transparency_texture[77][46] = 1;	doodle_left_transparency_texture[77][47] = 1;	doodle_left_transparency_texture[77][48] = 1;	doodle_left_transparency_texture[77][49] = 1;	doodle_left_transparency_texture[77][50] = 1;	doodle_left_transparency_texture[77][51] = 1;	doodle_left_transparency_texture[77][52] = 1;	doodle_left_transparency_texture[77][53] = 1;	doodle_left_transparency_texture[77][54] = 1;	doodle_left_transparency_texture[77][55] = 1;	doodle_left_transparency_texture[77][56] = 1;	doodle_left_transparency_texture[77][57] = 1;	doodle_left_transparency_texture[77][58] = 1;	doodle_left_transparency_texture[77][59] = 1;	doodle_left_transparency_texture[77][60] = 1;	doodle_left_transparency_texture[77][61] = 1;	doodle_left_transparency_texture[77][62] = 1;	doodle_left_transparency_texture[77][63] = 1;	doodle_left_transparency_texture[77][64] = 1;	doodle_left_transparency_texture[77][65] = 1;	doodle_left_transparency_texture[77][66] = 1;	doodle_left_transparency_texture[77][67] = 1;	doodle_left_transparency_texture[77][68] = 1;	doodle_left_transparency_texture[77][69] = 1;	doodle_left_transparency_texture[77][70] = 1;	doodle_left_transparency_texture[77][71] = 1;	doodle_left_transparency_texture[77][72] = 1;	doodle_left_transparency_texture[77][73] = 1;	doodle_left_transparency_texture[77][74] = 1;	doodle_left_transparency_texture[77][75] = 1;	doodle_left_transparency_texture[77][76] = 1;	doodle_left_transparency_texture[77][77] = 1;	doodle_left_transparency_texture[77][78] = 1;	doodle_left_transparency_texture[77][79] = 1;	doodle_left_transparency_texture[78][0] = 1;	doodle_left_transparency_texture[78][1] = 1;	doodle_left_transparency_texture[78][2] = 1;	doodle_left_transparency_texture[78][3] = 1;	doodle_left_transparency_texture[78][4] = 1;	doodle_left_transparency_texture[78][5] = 1;	doodle_left_transparency_texture[78][6] = 1;	doodle_left_transparency_texture[78][7] = 1;	doodle_left_transparency_texture[78][8] = 1;	doodle_left_transparency_texture[78][9] = 1;	doodle_left_transparency_texture[78][10] = 1;	doodle_left_transparency_texture[78][11] = 1;	doodle_left_transparency_texture[78][12] = 1;	doodle_left_transparency_texture[78][13] = 1;	doodle_left_transparency_texture[78][14] = 1;	doodle_left_transparency_texture[78][15] = 1;	doodle_left_transparency_texture[78][16] = 1;	doodle_left_transparency_texture[78][17] = 1;	doodle_left_transparency_texture[78][18] = 1;	doodle_left_transparency_texture[78][19] = 1;	doodle_left_transparency_texture[78][20] = 1;	doodle_left_transparency_texture[78][21] = 1;	doodle_left_transparency_texture[78][22] = 1;	doodle_left_transparency_texture[78][23] = 1;	doodle_left_transparency_texture[78][24] = 1;	doodle_left_transparency_texture[78][25] = 1;	doodle_left_transparency_texture[78][26] = 1;	doodle_left_transparency_texture[78][27] = 1;	doodle_left_transparency_texture[78][28] = 1;	doodle_left_transparency_texture[78][29] = 1;	doodle_left_transparency_texture[78][30] = 1;	doodle_left_transparency_texture[78][31] = 1;	doodle_left_transparency_texture[78][32] = 1;	doodle_left_transparency_texture[78][33] = 1;	doodle_left_transparency_texture[78][34] = 1;	doodle_left_transparency_texture[78][35] = 1;	doodle_left_transparency_texture[78][36] = 1;	doodle_left_transparency_texture[78][37] = 1;	doodle_left_transparency_texture[78][38] = 1;	doodle_left_transparency_texture[78][39] = 1;	doodle_left_transparency_texture[78][40] = 1;	doodle_left_transparency_texture[78][41] = 1;	doodle_left_transparency_texture[78][42] = 1;	doodle_left_transparency_texture[78][43] = 1;	doodle_left_transparency_texture[78][44] = 1;	doodle_left_transparency_texture[78][45] = 1;	doodle_left_transparency_texture[78][46] = 1;	doodle_left_transparency_texture[78][47] = 1;	doodle_left_transparency_texture[78][48] = 1;	doodle_left_transparency_texture[78][49] = 1;	doodle_left_transparency_texture[78][50] = 1;	doodle_left_transparency_texture[78][51] = 1;	doodle_left_transparency_texture[78][52] = 1;	doodle_left_transparency_texture[78][53] = 1;	doodle_left_transparency_texture[78][54] = 1;	doodle_left_transparency_texture[78][55] = 1;	doodle_left_transparency_texture[78][56] = 1;	doodle_left_transparency_texture[78][57] = 1;	doodle_left_transparency_texture[78][58] = 1;	doodle_left_transparency_texture[78][59] = 1;	doodle_left_transparency_texture[78][60] = 1;	doodle_left_transparency_texture[78][61] = 1;	doodle_left_transparency_texture[78][62] = 1;	doodle_left_transparency_texture[78][63] = 1;	doodle_left_transparency_texture[78][64] = 1;	doodle_left_transparency_texture[78][65] = 1;	doodle_left_transparency_texture[78][66] = 1;	doodle_left_transparency_texture[78][67] = 1;	doodle_left_transparency_texture[78][68] = 1;	doodle_left_transparency_texture[78][69] = 1;	doodle_left_transparency_texture[78][70] = 1;	doodle_left_transparency_texture[78][71] = 1;	doodle_left_transparency_texture[78][72] = 1;	doodle_left_transparency_texture[78][73] = 1;	doodle_left_transparency_texture[78][74] = 1;	doodle_left_transparency_texture[78][75] = 1;	doodle_left_transparency_texture[78][76] = 1;	doodle_left_transparency_texture[78][77] = 1;	doodle_left_transparency_texture[78][78] = 1;	doodle_left_transparency_texture[78][79] = 1;	doodle_left_transparency_texture[79][0] = 1;	doodle_left_transparency_texture[79][1] = 1;	doodle_left_transparency_texture[79][2] = 1;	doodle_left_transparency_texture[79][3] = 1;	doodle_left_transparency_texture[79][4] = 1;	doodle_left_transparency_texture[79][5] = 1;	doodle_left_transparency_texture[79][6] = 1;	doodle_left_transparency_texture[79][7] = 1;	doodle_left_transparency_texture[79][8] = 1;	doodle_left_transparency_texture[79][9] = 1;	doodle_left_transparency_texture[79][10] = 1;	doodle_left_transparency_texture[79][11] = 1;	doodle_left_transparency_texture[79][12] = 1;	doodle_left_transparency_texture[79][13] = 1;	doodle_left_transparency_texture[79][14] = 1;	doodle_left_transparency_texture[79][15] = 1;	doodle_left_transparency_texture[79][16] = 1;	doodle_left_transparency_texture[79][17] = 1;	doodle_left_transparency_texture[79][18] = 1;	doodle_left_transparency_texture[79][19] = 1;	doodle_left_transparency_texture[79][20] = 1;	doodle_left_transparency_texture[79][21] = 1;	doodle_left_transparency_texture[79][22] = 1;	doodle_left_transparency_texture[79][23] = 1;	doodle_left_transparency_texture[79][24] = 1;	doodle_left_transparency_texture[79][25] = 1;	doodle_left_transparency_texture[79][26] = 1;	doodle_left_transparency_texture[79][27] = 1;	doodle_left_transparency_texture[79][28] = 1;	doodle_left_transparency_texture[79][29] = 1;	doodle_left_transparency_texture[79][30] = 1;	doodle_left_transparency_texture[79][31] = 1;	doodle_left_transparency_texture[79][32] = 1;	doodle_left_transparency_texture[79][33] = 1;	doodle_left_transparency_texture[79][34] = 1;	doodle_left_transparency_texture[79][35] = 1;	doodle_left_transparency_texture[79][36] = 1;	doodle_left_transparency_texture[79][37] = 1;	doodle_left_transparency_texture[79][38] = 1;	doodle_left_transparency_texture[79][39] = 1;	doodle_left_transparency_texture[79][40] = 1;	doodle_left_transparency_texture[79][41] = 1;	doodle_left_transparency_texture[79][42] = 1;	doodle_left_transparency_texture[79][43] = 1;	doodle_left_transparency_texture[79][44] = 1;	doodle_left_transparency_texture[79][45] = 1;	doodle_left_transparency_texture[79][46] = 1;	doodle_left_transparency_texture[79][47] = 1;	doodle_left_transparency_texture[79][48] = 1;	doodle_left_transparency_texture[79][49] = 1;	doodle_left_transparency_texture[79][50] = 1;	doodle_left_transparency_texture[79][51] = 1;	doodle_left_transparency_texture[79][52] = 1;	doodle_left_transparency_texture[79][53] = 1;	doodle_left_transparency_texture[79][54] = 1;	doodle_left_transparency_texture[79][55] = 1;	doodle_left_transparency_texture[79][56] = 1;	doodle_left_transparency_texture[79][57] = 1;	doodle_left_transparency_texture[79][58] = 1;	doodle_left_transparency_texture[79][59] = 1;	doodle_left_transparency_texture[79][60] = 1;	doodle_left_transparency_texture[79][61] = 1;	doodle_left_transparency_texture[79][62] = 1;	doodle_left_transparency_texture[79][63] = 1;	doodle_left_transparency_texture[79][64] = 1;	doodle_left_transparency_texture[79][65] = 1;	doodle_left_transparency_texture[79][66] = 1;	doodle_left_transparency_texture[79][67] = 1;	doodle_left_transparency_texture[79][68] = 1;	doodle_left_transparency_texture[79][69] = 1;	doodle_left_transparency_texture[79][70] = 1;	doodle_left_transparency_texture[79][71] = 1;	doodle_left_transparency_texture[79][72] = 1;	doodle_left_transparency_texture[79][73] = 1;	doodle_left_transparency_texture[79][74] = 1;	doodle_left_transparency_texture[79][75] = 1;	doodle_left_transparency_texture[79][76] = 1;	doodle_left_transparency_texture[79][77] = 1;	doodle_left_transparency_texture[79][78] = 1;	doodle_left_transparency_texture[79][79] = 1;
end

endmodule