module signa(

);



endmodule
