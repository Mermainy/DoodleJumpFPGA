module board_specific(
	input MAX10_CLK1_50,
	
	output clk
);

assign clk = MAX10_CLK1_50;

endmodule
