`ifndef INITIAL_PLATFORM_GREEN

// Module definition:
// logic [29:0][99:0][2:0][3:0] platform_green_rgb;
// logic [29:0][99:0] platform_green_alpha;

`define INITIAL_PLATFORM_GREEN \
always_comb begin \
	platform_green_rgb[0][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[0][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[1][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[2][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[3][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[4][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[5][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[6][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[7][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[8][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[9][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[10][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[10][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[11][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[11][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[12][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[12][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[13][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[13][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[14][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[14][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[15][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[15][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[16][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[16][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[17][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[17][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[18][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[18][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][10] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][11] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][12] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][13] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][14] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][15] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][16] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][17] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][18] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][19] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][20] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][21] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][22] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][23] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][24] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][25] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][26] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][27] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][28] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][29] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][30] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][31] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][32] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][33] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][34] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][35] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][36] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][37] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][38] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][39] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][40] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][41] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][42] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][43] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][44] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][45] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][46] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][47] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][48] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][49] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][50] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][51] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][52] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][53] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][54] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][55] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][56] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][57] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][58] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][59] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][60] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][61] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][62] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][63] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][64] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][65] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][66] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][67] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][68] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][69] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][70] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][71] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][72] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][73] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][74] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][75] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][76] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][77] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][78] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][79] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][80] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][81] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][82] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][83] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][84] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][85] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][86] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][87] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][88] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][89] = {4'b0, 4'b1111, 4'b0}; \
	platform_green_rgb[19][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[19][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[20][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[21][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[22][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[23][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[24][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[25][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[26][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[27][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[28][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][0] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][1] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][2] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][3] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][4] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][5] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][6] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][7] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][8] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][9] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][10] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][11] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][12] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][13] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][14] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][15] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][16] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][17] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][18] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][19] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][20] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][21] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][22] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][23] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][24] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][25] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][26] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][27] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][28] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][29] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][30] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][31] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][32] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][33] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][34] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][35] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][36] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][37] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][38] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][39] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][40] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][41] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][42] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][43] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][44] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][45] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][46] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][47] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][48] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][49] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][50] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][51] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][52] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][53] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][54] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][55] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][56] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][57] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][58] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][59] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][60] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][61] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][62] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][63] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][64] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][65] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][66] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][67] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][68] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][69] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][70] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][71] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][72] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][73] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][74] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][75] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][76] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][77] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][78] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][79] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][80] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][81] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][82] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][83] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][84] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][85] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][86] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][87] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][88] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][89] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][90] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][91] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][92] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][93] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][94] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][95] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][96] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][97] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][98] = {4'b0, 4'b0, 4'b0}; \
	platform_green_rgb[29][99] = {4'b0, 4'b0, 4'b0}; \
	platform_green_alpha[0][0] = 1'b1; \
	platform_green_alpha[0][1] = 1'b1; \
	platform_green_alpha[0][2] = 1'b1; \
	platform_green_alpha[0][3] = 1'b1; \
	platform_green_alpha[0][4] = 1'b1; \
	platform_green_alpha[0][5] = 1'b1; \
	platform_green_alpha[0][6] = 1'b1; \
	platform_green_alpha[0][7] = 1'b1; \
	platform_green_alpha[0][8] = 1'b1; \
	platform_green_alpha[0][9] = 1'b1; \
	platform_green_alpha[0][10] = 1'b1; \
	platform_green_alpha[0][11] = 1'b1; \
	platform_green_alpha[0][12] = 1'b1; \
	platform_green_alpha[0][13] = 1'b1; \
	platform_green_alpha[0][14] = 1'b1; \
	platform_green_alpha[0][15] = 1'b1; \
	platform_green_alpha[0][16] = 1'b1; \
	platform_green_alpha[0][17] = 1'b1; \
	platform_green_alpha[0][18] = 1'b1; \
	platform_green_alpha[0][19] = 1'b1; \
	platform_green_alpha[0][20] = 1'b1; \
	platform_green_alpha[0][21] = 1'b1; \
	platform_green_alpha[0][22] = 1'b1; \
	platform_green_alpha[0][23] = 1'b1; \
	platform_green_alpha[0][24] = 1'b1; \
	platform_green_alpha[0][25] = 1'b1; \
	platform_green_alpha[0][26] = 1'b1; \
	platform_green_alpha[0][27] = 1'b1; \
	platform_green_alpha[0][28] = 1'b1; \
	platform_green_alpha[0][29] = 1'b1; \
	platform_green_alpha[0][30] = 1'b1; \
	platform_green_alpha[0][31] = 1'b1; \
	platform_green_alpha[0][32] = 1'b1; \
	platform_green_alpha[0][33] = 1'b1; \
	platform_green_alpha[0][34] = 1'b1; \
	platform_green_alpha[0][35] = 1'b1; \
	platform_green_alpha[0][36] = 1'b1; \
	platform_green_alpha[0][37] = 1'b1; \
	platform_green_alpha[0][38] = 1'b1; \
	platform_green_alpha[0][39] = 1'b1; \
	platform_green_alpha[0][40] = 1'b1; \
	platform_green_alpha[0][41] = 1'b1; \
	platform_green_alpha[0][42] = 1'b1; \
	platform_green_alpha[0][43] = 1'b1; \
	platform_green_alpha[0][44] = 1'b1; \
	platform_green_alpha[0][45] = 1'b1; \
	platform_green_alpha[0][46] = 1'b1; \
	platform_green_alpha[0][47] = 1'b1; \
	platform_green_alpha[0][48] = 1'b1; \
	platform_green_alpha[0][49] = 1'b1; \
	platform_green_alpha[0][50] = 1'b1; \
	platform_green_alpha[0][51] = 1'b1; \
	platform_green_alpha[0][52] = 1'b1; \
	platform_green_alpha[0][53] = 1'b1; \
	platform_green_alpha[0][54] = 1'b1; \
	platform_green_alpha[0][55] = 1'b1; \
	platform_green_alpha[0][56] = 1'b1; \
	platform_green_alpha[0][57] = 1'b1; \
	platform_green_alpha[0][58] = 1'b1; \
	platform_green_alpha[0][59] = 1'b1; \
	platform_green_alpha[0][60] = 1'b1; \
	platform_green_alpha[0][61] = 1'b1; \
	platform_green_alpha[0][62] = 1'b1; \
	platform_green_alpha[0][63] = 1'b1; \
	platform_green_alpha[0][64] = 1'b1; \
	platform_green_alpha[0][65] = 1'b1; \
	platform_green_alpha[0][66] = 1'b1; \
	platform_green_alpha[0][67] = 1'b1; \
	platform_green_alpha[0][68] = 1'b1; \
	platform_green_alpha[0][69] = 1'b1; \
	platform_green_alpha[0][70] = 1'b1; \
	platform_green_alpha[0][71] = 1'b1; \
	platform_green_alpha[0][72] = 1'b1; \
	platform_green_alpha[0][73] = 1'b1; \
	platform_green_alpha[0][74] = 1'b1; \
	platform_green_alpha[0][75] = 1'b1; \
	platform_green_alpha[0][76] = 1'b1; \
	platform_green_alpha[0][77] = 1'b1; \
	platform_green_alpha[0][78] = 1'b1; \
	platform_green_alpha[0][79] = 1'b1; \
	platform_green_alpha[0][80] = 1'b1; \
	platform_green_alpha[0][81] = 1'b1; \
	platform_green_alpha[0][82] = 1'b1; \
	platform_green_alpha[0][83] = 1'b1; \
	platform_green_alpha[0][84] = 1'b1; \
	platform_green_alpha[0][85] = 1'b1; \
	platform_green_alpha[0][86] = 1'b1; \
	platform_green_alpha[0][87] = 1'b1; \
	platform_green_alpha[0][88] = 1'b1; \
	platform_green_alpha[0][89] = 1'b1; \
	platform_green_alpha[0][90] = 1'b1; \
	platform_green_alpha[0][91] = 1'b1; \
	platform_green_alpha[0][92] = 1'b1; \
	platform_green_alpha[0][93] = 1'b1; \
	platform_green_alpha[0][94] = 1'b1; \
	platform_green_alpha[0][95] = 1'b1; \
	platform_green_alpha[0][96] = 1'b1; \
	platform_green_alpha[0][97] = 1'b1; \
	platform_green_alpha[0][98] = 1'b1; \
	platform_green_alpha[0][99] = 1'b1; \
	platform_green_alpha[1][0] = 1'b1; \
	platform_green_alpha[1][1] = 1'b1; \
	platform_green_alpha[1][2] = 1'b1; \
	platform_green_alpha[1][3] = 1'b1; \
	platform_green_alpha[1][4] = 1'b1; \
	platform_green_alpha[1][5] = 1'b1; \
	platform_green_alpha[1][6] = 1'b1; \
	platform_green_alpha[1][7] = 1'b1; \
	platform_green_alpha[1][8] = 1'b1; \
	platform_green_alpha[1][9] = 1'b1; \
	platform_green_alpha[1][10] = 1'b1; \
	platform_green_alpha[1][11] = 1'b1; \
	platform_green_alpha[1][12] = 1'b1; \
	platform_green_alpha[1][13] = 1'b1; \
	platform_green_alpha[1][14] = 1'b1; \
	platform_green_alpha[1][15] = 1'b1; \
	platform_green_alpha[1][16] = 1'b1; \
	platform_green_alpha[1][17] = 1'b1; \
	platform_green_alpha[1][18] = 1'b1; \
	platform_green_alpha[1][19] = 1'b1; \
	platform_green_alpha[1][20] = 1'b1; \
	platform_green_alpha[1][21] = 1'b1; \
	platform_green_alpha[1][22] = 1'b1; \
	platform_green_alpha[1][23] = 1'b1; \
	platform_green_alpha[1][24] = 1'b1; \
	platform_green_alpha[1][25] = 1'b1; \
	platform_green_alpha[1][26] = 1'b1; \
	platform_green_alpha[1][27] = 1'b1; \
	platform_green_alpha[1][28] = 1'b1; \
	platform_green_alpha[1][29] = 1'b1; \
	platform_green_alpha[1][30] = 1'b1; \
	platform_green_alpha[1][31] = 1'b1; \
	platform_green_alpha[1][32] = 1'b1; \
	platform_green_alpha[1][33] = 1'b1; \
	platform_green_alpha[1][34] = 1'b1; \
	platform_green_alpha[1][35] = 1'b1; \
	platform_green_alpha[1][36] = 1'b1; \
	platform_green_alpha[1][37] = 1'b1; \
	platform_green_alpha[1][38] = 1'b1; \
	platform_green_alpha[1][39] = 1'b1; \
	platform_green_alpha[1][40] = 1'b1; \
	platform_green_alpha[1][41] = 1'b1; \
	platform_green_alpha[1][42] = 1'b1; \
	platform_green_alpha[1][43] = 1'b1; \
	platform_green_alpha[1][44] = 1'b1; \
	platform_green_alpha[1][45] = 1'b1; \
	platform_green_alpha[1][46] = 1'b1; \
	platform_green_alpha[1][47] = 1'b1; \
	platform_green_alpha[1][48] = 1'b1; \
	platform_green_alpha[1][49] = 1'b1; \
	platform_green_alpha[1][50] = 1'b1; \
	platform_green_alpha[1][51] = 1'b1; \
	platform_green_alpha[1][52] = 1'b1; \
	platform_green_alpha[1][53] = 1'b1; \
	platform_green_alpha[1][54] = 1'b1; \
	platform_green_alpha[1][55] = 1'b1; \
	platform_green_alpha[1][56] = 1'b1; \
	platform_green_alpha[1][57] = 1'b1; \
	platform_green_alpha[1][58] = 1'b1; \
	platform_green_alpha[1][59] = 1'b1; \
	platform_green_alpha[1][60] = 1'b1; \
	platform_green_alpha[1][61] = 1'b1; \
	platform_green_alpha[1][62] = 1'b1; \
	platform_green_alpha[1][63] = 1'b1; \
	platform_green_alpha[1][64] = 1'b1; \
	platform_green_alpha[1][65] = 1'b1; \
	platform_green_alpha[1][66] = 1'b1; \
	platform_green_alpha[1][67] = 1'b1; \
	platform_green_alpha[1][68] = 1'b1; \
	platform_green_alpha[1][69] = 1'b1; \
	platform_green_alpha[1][70] = 1'b1; \
	platform_green_alpha[1][71] = 1'b1; \
	platform_green_alpha[1][72] = 1'b1; \
	platform_green_alpha[1][73] = 1'b1; \
	platform_green_alpha[1][74] = 1'b1; \
	platform_green_alpha[1][75] = 1'b1; \
	platform_green_alpha[1][76] = 1'b1; \
	platform_green_alpha[1][77] = 1'b1; \
	platform_green_alpha[1][78] = 1'b1; \
	platform_green_alpha[1][79] = 1'b1; \
	platform_green_alpha[1][80] = 1'b1; \
	platform_green_alpha[1][81] = 1'b1; \
	platform_green_alpha[1][82] = 1'b1; \
	platform_green_alpha[1][83] = 1'b1; \
	platform_green_alpha[1][84] = 1'b1; \
	platform_green_alpha[1][85] = 1'b1; \
	platform_green_alpha[1][86] = 1'b1; \
	platform_green_alpha[1][87] = 1'b1; \
	platform_green_alpha[1][88] = 1'b1; \
	platform_green_alpha[1][89] = 1'b1; \
	platform_green_alpha[1][90] = 1'b1; \
	platform_green_alpha[1][91] = 1'b1; \
	platform_green_alpha[1][92] = 1'b1; \
	platform_green_alpha[1][93] = 1'b1; \
	platform_green_alpha[1][94] = 1'b1; \
	platform_green_alpha[1][95] = 1'b1; \
	platform_green_alpha[1][96] = 1'b1; \
	platform_green_alpha[1][97] = 1'b1; \
	platform_green_alpha[1][98] = 1'b1; \
	platform_green_alpha[1][99] = 1'b1; \
	platform_green_alpha[2][0] = 1'b1; \
	platform_green_alpha[2][1] = 1'b1; \
	platform_green_alpha[2][2] = 1'b1; \
	platform_green_alpha[2][3] = 1'b1; \
	platform_green_alpha[2][4] = 1'b1; \
	platform_green_alpha[2][5] = 1'b1; \
	platform_green_alpha[2][6] = 1'b1; \
	platform_green_alpha[2][7] = 1'b1; \
	platform_green_alpha[2][8] = 1'b1; \
	platform_green_alpha[2][9] = 1'b1; \
	platform_green_alpha[2][10] = 1'b1; \
	platform_green_alpha[2][11] = 1'b1; \
	platform_green_alpha[2][12] = 1'b1; \
	platform_green_alpha[2][13] = 1'b1; \
	platform_green_alpha[2][14] = 1'b1; \
	platform_green_alpha[2][15] = 1'b1; \
	platform_green_alpha[2][16] = 1'b1; \
	platform_green_alpha[2][17] = 1'b1; \
	platform_green_alpha[2][18] = 1'b1; \
	platform_green_alpha[2][19] = 1'b1; \
	platform_green_alpha[2][20] = 1'b1; \
	platform_green_alpha[2][21] = 1'b1; \
	platform_green_alpha[2][22] = 1'b1; \
	platform_green_alpha[2][23] = 1'b1; \
	platform_green_alpha[2][24] = 1'b1; \
	platform_green_alpha[2][25] = 1'b1; \
	platform_green_alpha[2][26] = 1'b1; \
	platform_green_alpha[2][27] = 1'b1; \
	platform_green_alpha[2][28] = 1'b1; \
	platform_green_alpha[2][29] = 1'b1; \
	platform_green_alpha[2][30] = 1'b1; \
	platform_green_alpha[2][31] = 1'b1; \
	platform_green_alpha[2][32] = 1'b1; \
	platform_green_alpha[2][33] = 1'b1; \
	platform_green_alpha[2][34] = 1'b1; \
	platform_green_alpha[2][35] = 1'b1; \
	platform_green_alpha[2][36] = 1'b1; \
	platform_green_alpha[2][37] = 1'b1; \
	platform_green_alpha[2][38] = 1'b1; \
	platform_green_alpha[2][39] = 1'b1; \
	platform_green_alpha[2][40] = 1'b1; \
	platform_green_alpha[2][41] = 1'b1; \
	platform_green_alpha[2][42] = 1'b1; \
	platform_green_alpha[2][43] = 1'b1; \
	platform_green_alpha[2][44] = 1'b1; \
	platform_green_alpha[2][45] = 1'b1; \
	platform_green_alpha[2][46] = 1'b1; \
	platform_green_alpha[2][47] = 1'b1; \
	platform_green_alpha[2][48] = 1'b1; \
	platform_green_alpha[2][49] = 1'b1; \
	platform_green_alpha[2][50] = 1'b1; \
	platform_green_alpha[2][51] = 1'b1; \
	platform_green_alpha[2][52] = 1'b1; \
	platform_green_alpha[2][53] = 1'b1; \
	platform_green_alpha[2][54] = 1'b1; \
	platform_green_alpha[2][55] = 1'b1; \
	platform_green_alpha[2][56] = 1'b1; \
	platform_green_alpha[2][57] = 1'b1; \
	platform_green_alpha[2][58] = 1'b1; \
	platform_green_alpha[2][59] = 1'b1; \
	platform_green_alpha[2][60] = 1'b1; \
	platform_green_alpha[2][61] = 1'b1; \
	platform_green_alpha[2][62] = 1'b1; \
	platform_green_alpha[2][63] = 1'b1; \
	platform_green_alpha[2][64] = 1'b1; \
	platform_green_alpha[2][65] = 1'b1; \
	platform_green_alpha[2][66] = 1'b1; \
	platform_green_alpha[2][67] = 1'b1; \
	platform_green_alpha[2][68] = 1'b1; \
	platform_green_alpha[2][69] = 1'b1; \
	platform_green_alpha[2][70] = 1'b1; \
	platform_green_alpha[2][71] = 1'b1; \
	platform_green_alpha[2][72] = 1'b1; \
	platform_green_alpha[2][73] = 1'b1; \
	platform_green_alpha[2][74] = 1'b1; \
	platform_green_alpha[2][75] = 1'b1; \
	platform_green_alpha[2][76] = 1'b1; \
	platform_green_alpha[2][77] = 1'b1; \
	platform_green_alpha[2][78] = 1'b1; \
	platform_green_alpha[2][79] = 1'b1; \
	platform_green_alpha[2][80] = 1'b1; \
	platform_green_alpha[2][81] = 1'b1; \
	platform_green_alpha[2][82] = 1'b1; \
	platform_green_alpha[2][83] = 1'b1; \
	platform_green_alpha[2][84] = 1'b1; \
	platform_green_alpha[2][85] = 1'b1; \
	platform_green_alpha[2][86] = 1'b1; \
	platform_green_alpha[2][87] = 1'b1; \
	platform_green_alpha[2][88] = 1'b1; \
	platform_green_alpha[2][89] = 1'b1; \
	platform_green_alpha[2][90] = 1'b1; \
	platform_green_alpha[2][91] = 1'b1; \
	platform_green_alpha[2][92] = 1'b1; \
	platform_green_alpha[2][93] = 1'b1; \
	platform_green_alpha[2][94] = 1'b1; \
	platform_green_alpha[2][95] = 1'b1; \
	platform_green_alpha[2][96] = 1'b1; \
	platform_green_alpha[2][97] = 1'b1; \
	platform_green_alpha[2][98] = 1'b1; \
	platform_green_alpha[2][99] = 1'b1; \
	platform_green_alpha[3][0] = 1'b1; \
	platform_green_alpha[3][1] = 1'b1; \
	platform_green_alpha[3][2] = 1'b1; \
	platform_green_alpha[3][3] = 1'b1; \
	platform_green_alpha[3][4] = 1'b1; \
	platform_green_alpha[3][5] = 1'b1; \
	platform_green_alpha[3][6] = 1'b1; \
	platform_green_alpha[3][7] = 1'b1; \
	platform_green_alpha[3][8] = 1'b1; \
	platform_green_alpha[3][9] = 1'b1; \
	platform_green_alpha[3][10] = 1'b1; \
	platform_green_alpha[3][11] = 1'b1; \
	platform_green_alpha[3][12] = 1'b1; \
	platform_green_alpha[3][13] = 1'b1; \
	platform_green_alpha[3][14] = 1'b1; \
	platform_green_alpha[3][15] = 1'b1; \
	platform_green_alpha[3][16] = 1'b1; \
	platform_green_alpha[3][17] = 1'b1; \
	platform_green_alpha[3][18] = 1'b1; \
	platform_green_alpha[3][19] = 1'b1; \
	platform_green_alpha[3][20] = 1'b1; \
	platform_green_alpha[3][21] = 1'b1; \
	platform_green_alpha[3][22] = 1'b1; \
	platform_green_alpha[3][23] = 1'b1; \
	platform_green_alpha[3][24] = 1'b1; \
	platform_green_alpha[3][25] = 1'b1; \
	platform_green_alpha[3][26] = 1'b1; \
	platform_green_alpha[3][27] = 1'b1; \
	platform_green_alpha[3][28] = 1'b1; \
	platform_green_alpha[3][29] = 1'b1; \
	platform_green_alpha[3][30] = 1'b1; \
	platform_green_alpha[3][31] = 1'b1; \
	platform_green_alpha[3][32] = 1'b1; \
	platform_green_alpha[3][33] = 1'b1; \
	platform_green_alpha[3][34] = 1'b1; \
	platform_green_alpha[3][35] = 1'b1; \
	platform_green_alpha[3][36] = 1'b1; \
	platform_green_alpha[3][37] = 1'b1; \
	platform_green_alpha[3][38] = 1'b1; \
	platform_green_alpha[3][39] = 1'b1; \
	platform_green_alpha[3][40] = 1'b1; \
	platform_green_alpha[3][41] = 1'b1; \
	platform_green_alpha[3][42] = 1'b1; \
	platform_green_alpha[3][43] = 1'b1; \
	platform_green_alpha[3][44] = 1'b1; \
	platform_green_alpha[3][45] = 1'b1; \
	platform_green_alpha[3][46] = 1'b1; \
	platform_green_alpha[3][47] = 1'b1; \
	platform_green_alpha[3][48] = 1'b1; \
	platform_green_alpha[3][49] = 1'b1; \
	platform_green_alpha[3][50] = 1'b1; \
	platform_green_alpha[3][51] = 1'b1; \
	platform_green_alpha[3][52] = 1'b1; \
	platform_green_alpha[3][53] = 1'b1; \
	platform_green_alpha[3][54] = 1'b1; \
	platform_green_alpha[3][55] = 1'b1; \
	platform_green_alpha[3][56] = 1'b1; \
	platform_green_alpha[3][57] = 1'b1; \
	platform_green_alpha[3][58] = 1'b1; \
	platform_green_alpha[3][59] = 1'b1; \
	platform_green_alpha[3][60] = 1'b1; \
	platform_green_alpha[3][61] = 1'b1; \
	platform_green_alpha[3][62] = 1'b1; \
	platform_green_alpha[3][63] = 1'b1; \
	platform_green_alpha[3][64] = 1'b1; \
	platform_green_alpha[3][65] = 1'b1; \
	platform_green_alpha[3][66] = 1'b1; \
	platform_green_alpha[3][67] = 1'b1; \
	platform_green_alpha[3][68] = 1'b1; \
	platform_green_alpha[3][69] = 1'b1; \
	platform_green_alpha[3][70] = 1'b1; \
	platform_green_alpha[3][71] = 1'b1; \
	platform_green_alpha[3][72] = 1'b1; \
	platform_green_alpha[3][73] = 1'b1; \
	platform_green_alpha[3][74] = 1'b1; \
	platform_green_alpha[3][75] = 1'b1; \
	platform_green_alpha[3][76] = 1'b1; \
	platform_green_alpha[3][77] = 1'b1; \
	platform_green_alpha[3][78] = 1'b1; \
	platform_green_alpha[3][79] = 1'b1; \
	platform_green_alpha[3][80] = 1'b1; \
	platform_green_alpha[3][81] = 1'b1; \
	platform_green_alpha[3][82] = 1'b1; \
	platform_green_alpha[3][83] = 1'b1; \
	platform_green_alpha[3][84] = 1'b1; \
	platform_green_alpha[3][85] = 1'b1; \
	platform_green_alpha[3][86] = 1'b1; \
	platform_green_alpha[3][87] = 1'b1; \
	platform_green_alpha[3][88] = 1'b1; \
	platform_green_alpha[3][89] = 1'b1; \
	platform_green_alpha[3][90] = 1'b1; \
	platform_green_alpha[3][91] = 1'b1; \
	platform_green_alpha[3][92] = 1'b1; \
	platform_green_alpha[3][93] = 1'b1; \
	platform_green_alpha[3][94] = 1'b1; \
	platform_green_alpha[3][95] = 1'b1; \
	platform_green_alpha[3][96] = 1'b1; \
	platform_green_alpha[3][97] = 1'b1; \
	platform_green_alpha[3][98] = 1'b1; \
	platform_green_alpha[3][99] = 1'b1; \
	platform_green_alpha[4][0] = 1'b1; \
	platform_green_alpha[4][1] = 1'b1; \
	platform_green_alpha[4][2] = 1'b1; \
	platform_green_alpha[4][3] = 1'b1; \
	platform_green_alpha[4][4] = 1'b1; \
	platform_green_alpha[4][5] = 1'b1; \
	platform_green_alpha[4][6] = 1'b1; \
	platform_green_alpha[4][7] = 1'b1; \
	platform_green_alpha[4][8] = 1'b1; \
	platform_green_alpha[4][9] = 1'b1; \
	platform_green_alpha[4][10] = 1'b1; \
	platform_green_alpha[4][11] = 1'b1; \
	platform_green_alpha[4][12] = 1'b1; \
	platform_green_alpha[4][13] = 1'b1; \
	platform_green_alpha[4][14] = 1'b1; \
	platform_green_alpha[4][15] = 1'b1; \
	platform_green_alpha[4][16] = 1'b1; \
	platform_green_alpha[4][17] = 1'b1; \
	platform_green_alpha[4][18] = 1'b1; \
	platform_green_alpha[4][19] = 1'b1; \
	platform_green_alpha[4][20] = 1'b1; \
	platform_green_alpha[4][21] = 1'b1; \
	platform_green_alpha[4][22] = 1'b1; \
	platform_green_alpha[4][23] = 1'b1; \
	platform_green_alpha[4][24] = 1'b1; \
	platform_green_alpha[4][25] = 1'b1; \
	platform_green_alpha[4][26] = 1'b1; \
	platform_green_alpha[4][27] = 1'b1; \
	platform_green_alpha[4][28] = 1'b1; \
	platform_green_alpha[4][29] = 1'b1; \
	platform_green_alpha[4][30] = 1'b1; \
	platform_green_alpha[4][31] = 1'b1; \
	platform_green_alpha[4][32] = 1'b1; \
	platform_green_alpha[4][33] = 1'b1; \
	platform_green_alpha[4][34] = 1'b1; \
	platform_green_alpha[4][35] = 1'b1; \
	platform_green_alpha[4][36] = 1'b1; \
	platform_green_alpha[4][37] = 1'b1; \
	platform_green_alpha[4][38] = 1'b1; \
	platform_green_alpha[4][39] = 1'b1; \
	platform_green_alpha[4][40] = 1'b1; \
	platform_green_alpha[4][41] = 1'b1; \
	platform_green_alpha[4][42] = 1'b1; \
	platform_green_alpha[4][43] = 1'b1; \
	platform_green_alpha[4][44] = 1'b1; \
	platform_green_alpha[4][45] = 1'b1; \
	platform_green_alpha[4][46] = 1'b1; \
	platform_green_alpha[4][47] = 1'b1; \
	platform_green_alpha[4][48] = 1'b1; \
	platform_green_alpha[4][49] = 1'b1; \
	platform_green_alpha[4][50] = 1'b1; \
	platform_green_alpha[4][51] = 1'b1; \
	platform_green_alpha[4][52] = 1'b1; \
	platform_green_alpha[4][53] = 1'b1; \
	platform_green_alpha[4][54] = 1'b1; \
	platform_green_alpha[4][55] = 1'b1; \
	platform_green_alpha[4][56] = 1'b1; \
	platform_green_alpha[4][57] = 1'b1; \
	platform_green_alpha[4][58] = 1'b1; \
	platform_green_alpha[4][59] = 1'b1; \
	platform_green_alpha[4][60] = 1'b1; \
	platform_green_alpha[4][61] = 1'b1; \
	platform_green_alpha[4][62] = 1'b1; \
	platform_green_alpha[4][63] = 1'b1; \
	platform_green_alpha[4][64] = 1'b1; \
	platform_green_alpha[4][65] = 1'b1; \
	platform_green_alpha[4][66] = 1'b1; \
	platform_green_alpha[4][67] = 1'b1; \
	platform_green_alpha[4][68] = 1'b1; \
	platform_green_alpha[4][69] = 1'b1; \
	platform_green_alpha[4][70] = 1'b1; \
	platform_green_alpha[4][71] = 1'b1; \
	platform_green_alpha[4][72] = 1'b1; \
	platform_green_alpha[4][73] = 1'b1; \
	platform_green_alpha[4][74] = 1'b1; \
	platform_green_alpha[4][75] = 1'b1; \
	platform_green_alpha[4][76] = 1'b1; \
	platform_green_alpha[4][77] = 1'b1; \
	platform_green_alpha[4][78] = 1'b1; \
	platform_green_alpha[4][79] = 1'b1; \
	platform_green_alpha[4][80] = 1'b1; \
	platform_green_alpha[4][81] = 1'b1; \
	platform_green_alpha[4][82] = 1'b1; \
	platform_green_alpha[4][83] = 1'b1; \
	platform_green_alpha[4][84] = 1'b1; \
	platform_green_alpha[4][85] = 1'b1; \
	platform_green_alpha[4][86] = 1'b1; \
	platform_green_alpha[4][87] = 1'b1; \
	platform_green_alpha[4][88] = 1'b1; \
	platform_green_alpha[4][89] = 1'b1; \
	platform_green_alpha[4][90] = 1'b1; \
	platform_green_alpha[4][91] = 1'b1; \
	platform_green_alpha[4][92] = 1'b1; \
	platform_green_alpha[4][93] = 1'b1; \
	platform_green_alpha[4][94] = 1'b1; \
	platform_green_alpha[4][95] = 1'b1; \
	platform_green_alpha[4][96] = 1'b1; \
	platform_green_alpha[4][97] = 1'b1; \
	platform_green_alpha[4][98] = 1'b1; \
	platform_green_alpha[4][99] = 1'b1; \
	platform_green_alpha[5][0] = 1'b1; \
	platform_green_alpha[5][1] = 1'b1; \
	platform_green_alpha[5][2] = 1'b1; \
	platform_green_alpha[5][3] = 1'b1; \
	platform_green_alpha[5][4] = 1'b1; \
	platform_green_alpha[5][5] = 1'b1; \
	platform_green_alpha[5][6] = 1'b1; \
	platform_green_alpha[5][7] = 1'b1; \
	platform_green_alpha[5][8] = 1'b1; \
	platform_green_alpha[5][9] = 1'b1; \
	platform_green_alpha[5][10] = 1'b0; \
	platform_green_alpha[5][11] = 1'b0; \
	platform_green_alpha[5][12] = 1'b0; \
	platform_green_alpha[5][13] = 1'b0; \
	platform_green_alpha[5][14] = 1'b0; \
	platform_green_alpha[5][15] = 1'b0; \
	platform_green_alpha[5][16] = 1'b0; \
	platform_green_alpha[5][17] = 1'b0; \
	platform_green_alpha[5][18] = 1'b0; \
	platform_green_alpha[5][19] = 1'b0; \
	platform_green_alpha[5][20] = 1'b0; \
	platform_green_alpha[5][21] = 1'b0; \
	platform_green_alpha[5][22] = 1'b0; \
	platform_green_alpha[5][23] = 1'b0; \
	platform_green_alpha[5][24] = 1'b0; \
	platform_green_alpha[5][25] = 1'b0; \
	platform_green_alpha[5][26] = 1'b0; \
	platform_green_alpha[5][27] = 1'b0; \
	platform_green_alpha[5][28] = 1'b0; \
	platform_green_alpha[5][29] = 1'b0; \
	platform_green_alpha[5][30] = 1'b0; \
	platform_green_alpha[5][31] = 1'b0; \
	platform_green_alpha[5][32] = 1'b0; \
	platform_green_alpha[5][33] = 1'b0; \
	platform_green_alpha[5][34] = 1'b0; \
	platform_green_alpha[5][35] = 1'b0; \
	platform_green_alpha[5][36] = 1'b0; \
	platform_green_alpha[5][37] = 1'b0; \
	platform_green_alpha[5][38] = 1'b0; \
	platform_green_alpha[5][39] = 1'b0; \
	platform_green_alpha[5][40] = 1'b0; \
	platform_green_alpha[5][41] = 1'b0; \
	platform_green_alpha[5][42] = 1'b0; \
	platform_green_alpha[5][43] = 1'b0; \
	platform_green_alpha[5][44] = 1'b0; \
	platform_green_alpha[5][45] = 1'b0; \
	platform_green_alpha[5][46] = 1'b0; \
	platform_green_alpha[5][47] = 1'b0; \
	platform_green_alpha[5][48] = 1'b0; \
	platform_green_alpha[5][49] = 1'b0; \
	platform_green_alpha[5][50] = 1'b0; \
	platform_green_alpha[5][51] = 1'b0; \
	platform_green_alpha[5][52] = 1'b0; \
	platform_green_alpha[5][53] = 1'b0; \
	platform_green_alpha[5][54] = 1'b0; \
	platform_green_alpha[5][55] = 1'b0; \
	platform_green_alpha[5][56] = 1'b0; \
	platform_green_alpha[5][57] = 1'b0; \
	platform_green_alpha[5][58] = 1'b0; \
	platform_green_alpha[5][59] = 1'b0; \
	platform_green_alpha[5][60] = 1'b0; \
	platform_green_alpha[5][61] = 1'b0; \
	platform_green_alpha[5][62] = 1'b0; \
	platform_green_alpha[5][63] = 1'b0; \
	platform_green_alpha[5][64] = 1'b0; \
	platform_green_alpha[5][65] = 1'b0; \
	platform_green_alpha[5][66] = 1'b0; \
	platform_green_alpha[5][67] = 1'b0; \
	platform_green_alpha[5][68] = 1'b0; \
	platform_green_alpha[5][69] = 1'b0; \
	platform_green_alpha[5][70] = 1'b0; \
	platform_green_alpha[5][71] = 1'b0; \
	platform_green_alpha[5][72] = 1'b0; \
	platform_green_alpha[5][73] = 1'b0; \
	platform_green_alpha[5][74] = 1'b0; \
	platform_green_alpha[5][75] = 1'b0; \
	platform_green_alpha[5][76] = 1'b0; \
	platform_green_alpha[5][77] = 1'b0; \
	platform_green_alpha[5][78] = 1'b0; \
	platform_green_alpha[5][79] = 1'b0; \
	platform_green_alpha[5][80] = 1'b0; \
	platform_green_alpha[5][81] = 1'b0; \
	platform_green_alpha[5][82] = 1'b0; \
	platform_green_alpha[5][83] = 1'b0; \
	platform_green_alpha[5][84] = 1'b0; \
	platform_green_alpha[5][85] = 1'b0; \
	platform_green_alpha[5][86] = 1'b0; \
	platform_green_alpha[5][87] = 1'b0; \
	platform_green_alpha[5][88] = 1'b0; \
	platform_green_alpha[5][89] = 1'b0; \
	platform_green_alpha[5][90] = 1'b1; \
	platform_green_alpha[5][91] = 1'b1; \
	platform_green_alpha[5][92] = 1'b1; \
	platform_green_alpha[5][93] = 1'b1; \
	platform_green_alpha[5][94] = 1'b1; \
	platform_green_alpha[5][95] = 1'b1; \
	platform_green_alpha[5][96] = 1'b1; \
	platform_green_alpha[5][97] = 1'b1; \
	platform_green_alpha[5][98] = 1'b1; \
	platform_green_alpha[5][99] = 1'b1; \
	platform_green_alpha[6][0] = 1'b1; \
	platform_green_alpha[6][1] = 1'b1; \
	platform_green_alpha[6][2] = 1'b1; \
	platform_green_alpha[6][3] = 1'b1; \
	platform_green_alpha[6][4] = 1'b1; \
	platform_green_alpha[6][5] = 1'b1; \
	platform_green_alpha[6][6] = 1'b1; \
	platform_green_alpha[6][7] = 1'b1; \
	platform_green_alpha[6][8] = 1'b1; \
	platform_green_alpha[6][9] = 1'b1; \
	platform_green_alpha[6][10] = 1'b0; \
	platform_green_alpha[6][11] = 1'b0; \
	platform_green_alpha[6][12] = 1'b0; \
	platform_green_alpha[6][13] = 1'b0; \
	platform_green_alpha[6][14] = 1'b0; \
	platform_green_alpha[6][15] = 1'b0; \
	platform_green_alpha[6][16] = 1'b0; \
	platform_green_alpha[6][17] = 1'b0; \
	platform_green_alpha[6][18] = 1'b0; \
	platform_green_alpha[6][19] = 1'b0; \
	platform_green_alpha[6][20] = 1'b0; \
	platform_green_alpha[6][21] = 1'b0; \
	platform_green_alpha[6][22] = 1'b0; \
	platform_green_alpha[6][23] = 1'b0; \
	platform_green_alpha[6][24] = 1'b0; \
	platform_green_alpha[6][25] = 1'b0; \
	platform_green_alpha[6][26] = 1'b0; \
	platform_green_alpha[6][27] = 1'b0; \
	platform_green_alpha[6][28] = 1'b0; \
	platform_green_alpha[6][29] = 1'b0; \
	platform_green_alpha[6][30] = 1'b0; \
	platform_green_alpha[6][31] = 1'b0; \
	platform_green_alpha[6][32] = 1'b0; \
	platform_green_alpha[6][33] = 1'b0; \
	platform_green_alpha[6][34] = 1'b0; \
	platform_green_alpha[6][35] = 1'b0; \
	platform_green_alpha[6][36] = 1'b0; \
	platform_green_alpha[6][37] = 1'b0; \
	platform_green_alpha[6][38] = 1'b0; \
	platform_green_alpha[6][39] = 1'b0; \
	platform_green_alpha[6][40] = 1'b0; \
	platform_green_alpha[6][41] = 1'b0; \
	platform_green_alpha[6][42] = 1'b0; \
	platform_green_alpha[6][43] = 1'b0; \
	platform_green_alpha[6][44] = 1'b0; \
	platform_green_alpha[6][45] = 1'b0; \
	platform_green_alpha[6][46] = 1'b0; \
	platform_green_alpha[6][47] = 1'b0; \
	platform_green_alpha[6][48] = 1'b0; \
	platform_green_alpha[6][49] = 1'b0; \
	platform_green_alpha[6][50] = 1'b0; \
	platform_green_alpha[6][51] = 1'b0; \
	platform_green_alpha[6][52] = 1'b0; \
	platform_green_alpha[6][53] = 1'b0; \
	platform_green_alpha[6][54] = 1'b0; \
	platform_green_alpha[6][55] = 1'b0; \
	platform_green_alpha[6][56] = 1'b0; \
	platform_green_alpha[6][57] = 1'b0; \
	platform_green_alpha[6][58] = 1'b0; \
	platform_green_alpha[6][59] = 1'b0; \
	platform_green_alpha[6][60] = 1'b0; \
	platform_green_alpha[6][61] = 1'b0; \
	platform_green_alpha[6][62] = 1'b0; \
	platform_green_alpha[6][63] = 1'b0; \
	platform_green_alpha[6][64] = 1'b0; \
	platform_green_alpha[6][65] = 1'b0; \
	platform_green_alpha[6][66] = 1'b0; \
	platform_green_alpha[6][67] = 1'b0; \
	platform_green_alpha[6][68] = 1'b0; \
	platform_green_alpha[6][69] = 1'b0; \
	platform_green_alpha[6][70] = 1'b0; \
	platform_green_alpha[6][71] = 1'b0; \
	platform_green_alpha[6][72] = 1'b0; \
	platform_green_alpha[6][73] = 1'b0; \
	platform_green_alpha[6][74] = 1'b0; \
	platform_green_alpha[6][75] = 1'b0; \
	platform_green_alpha[6][76] = 1'b0; \
	platform_green_alpha[6][77] = 1'b0; \
	platform_green_alpha[6][78] = 1'b0; \
	platform_green_alpha[6][79] = 1'b0; \
	platform_green_alpha[6][80] = 1'b0; \
	platform_green_alpha[6][81] = 1'b0; \
	platform_green_alpha[6][82] = 1'b0; \
	platform_green_alpha[6][83] = 1'b0; \
	platform_green_alpha[6][84] = 1'b0; \
	platform_green_alpha[6][85] = 1'b0; \
	platform_green_alpha[6][86] = 1'b0; \
	platform_green_alpha[6][87] = 1'b0; \
	platform_green_alpha[6][88] = 1'b0; \
	platform_green_alpha[6][89] = 1'b0; \
	platform_green_alpha[6][90] = 1'b1; \
	platform_green_alpha[6][91] = 1'b1; \
	platform_green_alpha[6][92] = 1'b1; \
	platform_green_alpha[6][93] = 1'b1; \
	platform_green_alpha[6][94] = 1'b1; \
	platform_green_alpha[6][95] = 1'b1; \
	platform_green_alpha[6][96] = 1'b1; \
	platform_green_alpha[6][97] = 1'b1; \
	platform_green_alpha[6][98] = 1'b1; \
	platform_green_alpha[6][99] = 1'b1; \
	platform_green_alpha[7][0] = 1'b1; \
	platform_green_alpha[7][1] = 1'b1; \
	platform_green_alpha[7][2] = 1'b1; \
	platform_green_alpha[7][3] = 1'b1; \
	platform_green_alpha[7][4] = 1'b1; \
	platform_green_alpha[7][5] = 1'b1; \
	platform_green_alpha[7][6] = 1'b1; \
	platform_green_alpha[7][7] = 1'b1; \
	platform_green_alpha[7][8] = 1'b1; \
	platform_green_alpha[7][9] = 1'b1; \
	platform_green_alpha[7][10] = 1'b0; \
	platform_green_alpha[7][11] = 1'b0; \
	platform_green_alpha[7][12] = 1'b0; \
	platform_green_alpha[7][13] = 1'b0; \
	platform_green_alpha[7][14] = 1'b0; \
	platform_green_alpha[7][15] = 1'b0; \
	platform_green_alpha[7][16] = 1'b0; \
	platform_green_alpha[7][17] = 1'b0; \
	platform_green_alpha[7][18] = 1'b0; \
	platform_green_alpha[7][19] = 1'b0; \
	platform_green_alpha[7][20] = 1'b0; \
	platform_green_alpha[7][21] = 1'b0; \
	platform_green_alpha[7][22] = 1'b0; \
	platform_green_alpha[7][23] = 1'b0; \
	platform_green_alpha[7][24] = 1'b0; \
	platform_green_alpha[7][25] = 1'b0; \
	platform_green_alpha[7][26] = 1'b0; \
	platform_green_alpha[7][27] = 1'b0; \
	platform_green_alpha[7][28] = 1'b0; \
	platform_green_alpha[7][29] = 1'b0; \
	platform_green_alpha[7][30] = 1'b0; \
	platform_green_alpha[7][31] = 1'b0; \
	platform_green_alpha[7][32] = 1'b0; \
	platform_green_alpha[7][33] = 1'b0; \
	platform_green_alpha[7][34] = 1'b0; \
	platform_green_alpha[7][35] = 1'b0; \
	platform_green_alpha[7][36] = 1'b0; \
	platform_green_alpha[7][37] = 1'b0; \
	platform_green_alpha[7][38] = 1'b0; \
	platform_green_alpha[7][39] = 1'b0; \
	platform_green_alpha[7][40] = 1'b0; \
	platform_green_alpha[7][41] = 1'b0; \
	platform_green_alpha[7][42] = 1'b0; \
	platform_green_alpha[7][43] = 1'b0; \
	platform_green_alpha[7][44] = 1'b0; \
	platform_green_alpha[7][45] = 1'b0; \
	platform_green_alpha[7][46] = 1'b0; \
	platform_green_alpha[7][47] = 1'b0; \
	platform_green_alpha[7][48] = 1'b0; \
	platform_green_alpha[7][49] = 1'b0; \
	platform_green_alpha[7][50] = 1'b0; \
	platform_green_alpha[7][51] = 1'b0; \
	platform_green_alpha[7][52] = 1'b0; \
	platform_green_alpha[7][53] = 1'b0; \
	platform_green_alpha[7][54] = 1'b0; \
	platform_green_alpha[7][55] = 1'b0; \
	platform_green_alpha[7][56] = 1'b0; \
	platform_green_alpha[7][57] = 1'b0; \
	platform_green_alpha[7][58] = 1'b0; \
	platform_green_alpha[7][59] = 1'b0; \
	platform_green_alpha[7][60] = 1'b0; \
	platform_green_alpha[7][61] = 1'b0; \
	platform_green_alpha[7][62] = 1'b0; \
	platform_green_alpha[7][63] = 1'b0; \
	platform_green_alpha[7][64] = 1'b0; \
	platform_green_alpha[7][65] = 1'b0; \
	platform_green_alpha[7][66] = 1'b0; \
	platform_green_alpha[7][67] = 1'b0; \
	platform_green_alpha[7][68] = 1'b0; \
	platform_green_alpha[7][69] = 1'b0; \
	platform_green_alpha[7][70] = 1'b0; \
	platform_green_alpha[7][71] = 1'b0; \
	platform_green_alpha[7][72] = 1'b0; \
	platform_green_alpha[7][73] = 1'b0; \
	platform_green_alpha[7][74] = 1'b0; \
	platform_green_alpha[7][75] = 1'b0; \
	platform_green_alpha[7][76] = 1'b0; \
	platform_green_alpha[7][77] = 1'b0; \
	platform_green_alpha[7][78] = 1'b0; \
	platform_green_alpha[7][79] = 1'b0; \
	platform_green_alpha[7][80] = 1'b0; \
	platform_green_alpha[7][81] = 1'b0; \
	platform_green_alpha[7][82] = 1'b0; \
	platform_green_alpha[7][83] = 1'b0; \
	platform_green_alpha[7][84] = 1'b0; \
	platform_green_alpha[7][85] = 1'b0; \
	platform_green_alpha[7][86] = 1'b0; \
	platform_green_alpha[7][87] = 1'b0; \
	platform_green_alpha[7][88] = 1'b0; \
	platform_green_alpha[7][89] = 1'b0; \
	platform_green_alpha[7][90] = 1'b1; \
	platform_green_alpha[7][91] = 1'b1; \
	platform_green_alpha[7][92] = 1'b1; \
	platform_green_alpha[7][93] = 1'b1; \
	platform_green_alpha[7][94] = 1'b1; \
	platform_green_alpha[7][95] = 1'b1; \
	platform_green_alpha[7][96] = 1'b1; \
	platform_green_alpha[7][97] = 1'b1; \
	platform_green_alpha[7][98] = 1'b1; \
	platform_green_alpha[7][99] = 1'b1; \
	platform_green_alpha[8][0] = 1'b1; \
	platform_green_alpha[8][1] = 1'b1; \
	platform_green_alpha[8][2] = 1'b1; \
	platform_green_alpha[8][3] = 1'b1; \
	platform_green_alpha[8][4] = 1'b1; \
	platform_green_alpha[8][5] = 1'b1; \
	platform_green_alpha[8][6] = 1'b1; \
	platform_green_alpha[8][7] = 1'b1; \
	platform_green_alpha[8][8] = 1'b1; \
	platform_green_alpha[8][9] = 1'b1; \
	platform_green_alpha[8][10] = 1'b0; \
	platform_green_alpha[8][11] = 1'b0; \
	platform_green_alpha[8][12] = 1'b0; \
	platform_green_alpha[8][13] = 1'b0; \
	platform_green_alpha[8][14] = 1'b0; \
	platform_green_alpha[8][15] = 1'b0; \
	platform_green_alpha[8][16] = 1'b0; \
	platform_green_alpha[8][17] = 1'b0; \
	platform_green_alpha[8][18] = 1'b0; \
	platform_green_alpha[8][19] = 1'b0; \
	platform_green_alpha[8][20] = 1'b0; \
	platform_green_alpha[8][21] = 1'b0; \
	platform_green_alpha[8][22] = 1'b0; \
	platform_green_alpha[8][23] = 1'b0; \
	platform_green_alpha[8][24] = 1'b0; \
	platform_green_alpha[8][25] = 1'b0; \
	platform_green_alpha[8][26] = 1'b0; \
	platform_green_alpha[8][27] = 1'b0; \
	platform_green_alpha[8][28] = 1'b0; \
	platform_green_alpha[8][29] = 1'b0; \
	platform_green_alpha[8][30] = 1'b0; \
	platform_green_alpha[8][31] = 1'b0; \
	platform_green_alpha[8][32] = 1'b0; \
	platform_green_alpha[8][33] = 1'b0; \
	platform_green_alpha[8][34] = 1'b0; \
	platform_green_alpha[8][35] = 1'b0; \
	platform_green_alpha[8][36] = 1'b0; \
	platform_green_alpha[8][37] = 1'b0; \
	platform_green_alpha[8][38] = 1'b0; \
	platform_green_alpha[8][39] = 1'b0; \
	platform_green_alpha[8][40] = 1'b0; \
	platform_green_alpha[8][41] = 1'b0; \
	platform_green_alpha[8][42] = 1'b0; \
	platform_green_alpha[8][43] = 1'b0; \
	platform_green_alpha[8][44] = 1'b0; \
	platform_green_alpha[8][45] = 1'b0; \
	platform_green_alpha[8][46] = 1'b0; \
	platform_green_alpha[8][47] = 1'b0; \
	platform_green_alpha[8][48] = 1'b0; \
	platform_green_alpha[8][49] = 1'b0; \
	platform_green_alpha[8][50] = 1'b0; \
	platform_green_alpha[8][51] = 1'b0; \
	platform_green_alpha[8][52] = 1'b0; \
	platform_green_alpha[8][53] = 1'b0; \
	platform_green_alpha[8][54] = 1'b0; \
	platform_green_alpha[8][55] = 1'b0; \
	platform_green_alpha[8][56] = 1'b0; \
	platform_green_alpha[8][57] = 1'b0; \
	platform_green_alpha[8][58] = 1'b0; \
	platform_green_alpha[8][59] = 1'b0; \
	platform_green_alpha[8][60] = 1'b0; \
	platform_green_alpha[8][61] = 1'b0; \
	platform_green_alpha[8][62] = 1'b0; \
	platform_green_alpha[8][63] = 1'b0; \
	platform_green_alpha[8][64] = 1'b0; \
	platform_green_alpha[8][65] = 1'b0; \
	platform_green_alpha[8][66] = 1'b0; \
	platform_green_alpha[8][67] = 1'b0; \
	platform_green_alpha[8][68] = 1'b0; \
	platform_green_alpha[8][69] = 1'b0; \
	platform_green_alpha[8][70] = 1'b0; \
	platform_green_alpha[8][71] = 1'b0; \
	platform_green_alpha[8][72] = 1'b0; \
	platform_green_alpha[8][73] = 1'b0; \
	platform_green_alpha[8][74] = 1'b0; \
	platform_green_alpha[8][75] = 1'b0; \
	platform_green_alpha[8][76] = 1'b0; \
	platform_green_alpha[8][77] = 1'b0; \
	platform_green_alpha[8][78] = 1'b0; \
	platform_green_alpha[8][79] = 1'b0; \
	platform_green_alpha[8][80] = 1'b0; \
	platform_green_alpha[8][81] = 1'b0; \
	platform_green_alpha[8][82] = 1'b0; \
	platform_green_alpha[8][83] = 1'b0; \
	platform_green_alpha[8][84] = 1'b0; \
	platform_green_alpha[8][85] = 1'b0; \
	platform_green_alpha[8][86] = 1'b0; \
	platform_green_alpha[8][87] = 1'b0; \
	platform_green_alpha[8][88] = 1'b0; \
	platform_green_alpha[8][89] = 1'b0; \
	platform_green_alpha[8][90] = 1'b1; \
	platform_green_alpha[8][91] = 1'b1; \
	platform_green_alpha[8][92] = 1'b1; \
	platform_green_alpha[8][93] = 1'b1; \
	platform_green_alpha[8][94] = 1'b1; \
	platform_green_alpha[8][95] = 1'b1; \
	platform_green_alpha[8][96] = 1'b1; \
	platform_green_alpha[8][97] = 1'b1; \
	platform_green_alpha[8][98] = 1'b1; \
	platform_green_alpha[8][99] = 1'b1; \
	platform_green_alpha[9][0] = 1'b1; \
	platform_green_alpha[9][1] = 1'b1; \
	platform_green_alpha[9][2] = 1'b1; \
	platform_green_alpha[9][3] = 1'b1; \
	platform_green_alpha[9][4] = 1'b1; \
	platform_green_alpha[9][5] = 1'b1; \
	platform_green_alpha[9][6] = 1'b1; \
	platform_green_alpha[9][7] = 1'b1; \
	platform_green_alpha[9][8] = 1'b1; \
	platform_green_alpha[9][9] = 1'b1; \
	platform_green_alpha[9][10] = 1'b0; \
	platform_green_alpha[9][11] = 1'b0; \
	platform_green_alpha[9][12] = 1'b0; \
	platform_green_alpha[9][13] = 1'b0; \
	platform_green_alpha[9][14] = 1'b0; \
	platform_green_alpha[9][15] = 1'b0; \
	platform_green_alpha[9][16] = 1'b0; \
	platform_green_alpha[9][17] = 1'b0; \
	platform_green_alpha[9][18] = 1'b0; \
	platform_green_alpha[9][19] = 1'b0; \
	platform_green_alpha[9][20] = 1'b0; \
	platform_green_alpha[9][21] = 1'b0; \
	platform_green_alpha[9][22] = 1'b0; \
	platform_green_alpha[9][23] = 1'b0; \
	platform_green_alpha[9][24] = 1'b0; \
	platform_green_alpha[9][25] = 1'b0; \
	platform_green_alpha[9][26] = 1'b0; \
	platform_green_alpha[9][27] = 1'b0; \
	platform_green_alpha[9][28] = 1'b0; \
	platform_green_alpha[9][29] = 1'b0; \
	platform_green_alpha[9][30] = 1'b0; \
	platform_green_alpha[9][31] = 1'b0; \
	platform_green_alpha[9][32] = 1'b0; \
	platform_green_alpha[9][33] = 1'b0; \
	platform_green_alpha[9][34] = 1'b0; \
	platform_green_alpha[9][35] = 1'b0; \
	platform_green_alpha[9][36] = 1'b0; \
	platform_green_alpha[9][37] = 1'b0; \
	platform_green_alpha[9][38] = 1'b0; \
	platform_green_alpha[9][39] = 1'b0; \
	platform_green_alpha[9][40] = 1'b0; \
	platform_green_alpha[9][41] = 1'b0; \
	platform_green_alpha[9][42] = 1'b0; \
	platform_green_alpha[9][43] = 1'b0; \
	platform_green_alpha[9][44] = 1'b0; \
	platform_green_alpha[9][45] = 1'b0; \
	platform_green_alpha[9][46] = 1'b0; \
	platform_green_alpha[9][47] = 1'b0; \
	platform_green_alpha[9][48] = 1'b0; \
	platform_green_alpha[9][49] = 1'b0; \
	platform_green_alpha[9][50] = 1'b0; \
	platform_green_alpha[9][51] = 1'b0; \
	platform_green_alpha[9][52] = 1'b0; \
	platform_green_alpha[9][53] = 1'b0; \
	platform_green_alpha[9][54] = 1'b0; \
	platform_green_alpha[9][55] = 1'b0; \
	platform_green_alpha[9][56] = 1'b0; \
	platform_green_alpha[9][57] = 1'b0; \
	platform_green_alpha[9][58] = 1'b0; \
	platform_green_alpha[9][59] = 1'b0; \
	platform_green_alpha[9][60] = 1'b0; \
	platform_green_alpha[9][61] = 1'b0; \
	platform_green_alpha[9][62] = 1'b0; \
	platform_green_alpha[9][63] = 1'b0; \
	platform_green_alpha[9][64] = 1'b0; \
	platform_green_alpha[9][65] = 1'b0; \
	platform_green_alpha[9][66] = 1'b0; \
	platform_green_alpha[9][67] = 1'b0; \
	platform_green_alpha[9][68] = 1'b0; \
	platform_green_alpha[9][69] = 1'b0; \
	platform_green_alpha[9][70] = 1'b0; \
	platform_green_alpha[9][71] = 1'b0; \
	platform_green_alpha[9][72] = 1'b0; \
	platform_green_alpha[9][73] = 1'b0; \
	platform_green_alpha[9][74] = 1'b0; \
	platform_green_alpha[9][75] = 1'b0; \
	platform_green_alpha[9][76] = 1'b0; \
	platform_green_alpha[9][77] = 1'b0; \
	platform_green_alpha[9][78] = 1'b0; \
	platform_green_alpha[9][79] = 1'b0; \
	platform_green_alpha[9][80] = 1'b0; \
	platform_green_alpha[9][81] = 1'b0; \
	platform_green_alpha[9][82] = 1'b0; \
	platform_green_alpha[9][83] = 1'b0; \
	platform_green_alpha[9][84] = 1'b0; \
	platform_green_alpha[9][85] = 1'b0; \
	platform_green_alpha[9][86] = 1'b0; \
	platform_green_alpha[9][87] = 1'b0; \
	platform_green_alpha[9][88] = 1'b0; \
	platform_green_alpha[9][89] = 1'b0; \
	platform_green_alpha[9][90] = 1'b1; \
	platform_green_alpha[9][91] = 1'b1; \
	platform_green_alpha[9][92] = 1'b1; \
	platform_green_alpha[9][93] = 1'b1; \
	platform_green_alpha[9][94] = 1'b1; \
	platform_green_alpha[9][95] = 1'b1; \
	platform_green_alpha[9][96] = 1'b1; \
	platform_green_alpha[9][97] = 1'b1; \
	platform_green_alpha[9][98] = 1'b1; \
	platform_green_alpha[9][99] = 1'b1; \
	platform_green_alpha[10][0] = 1'b1; \
	platform_green_alpha[10][1] = 1'b1; \
	platform_green_alpha[10][2] = 1'b1; \
	platform_green_alpha[10][3] = 1'b1; \
	platform_green_alpha[10][4] = 1'b1; \
	platform_green_alpha[10][5] = 1'b0; \
	platform_green_alpha[10][6] = 1'b0; \
	platform_green_alpha[10][7] = 1'b0; \
	platform_green_alpha[10][8] = 1'b0; \
	platform_green_alpha[10][9] = 1'b0; \
	platform_green_alpha[10][10] = 1'b0; \
	platform_green_alpha[10][11] = 1'b0; \
	platform_green_alpha[10][12] = 1'b0; \
	platform_green_alpha[10][13] = 1'b0; \
	platform_green_alpha[10][14] = 1'b0; \
	platform_green_alpha[10][15] = 1'b0; \
	platform_green_alpha[10][16] = 1'b0; \
	platform_green_alpha[10][17] = 1'b0; \
	platform_green_alpha[10][18] = 1'b0; \
	platform_green_alpha[10][19] = 1'b0; \
	platform_green_alpha[10][20] = 1'b0; \
	platform_green_alpha[10][21] = 1'b0; \
	platform_green_alpha[10][22] = 1'b0; \
	platform_green_alpha[10][23] = 1'b0; \
	platform_green_alpha[10][24] = 1'b0; \
	platform_green_alpha[10][25] = 1'b0; \
	platform_green_alpha[10][26] = 1'b0; \
	platform_green_alpha[10][27] = 1'b0; \
	platform_green_alpha[10][28] = 1'b0; \
	platform_green_alpha[10][29] = 1'b0; \
	platform_green_alpha[10][30] = 1'b0; \
	platform_green_alpha[10][31] = 1'b0; \
	platform_green_alpha[10][32] = 1'b0; \
	platform_green_alpha[10][33] = 1'b0; \
	platform_green_alpha[10][34] = 1'b0; \
	platform_green_alpha[10][35] = 1'b0; \
	platform_green_alpha[10][36] = 1'b0; \
	platform_green_alpha[10][37] = 1'b0; \
	platform_green_alpha[10][38] = 1'b0; \
	platform_green_alpha[10][39] = 1'b0; \
	platform_green_alpha[10][40] = 1'b0; \
	platform_green_alpha[10][41] = 1'b0; \
	platform_green_alpha[10][42] = 1'b0; \
	platform_green_alpha[10][43] = 1'b0; \
	platform_green_alpha[10][44] = 1'b0; \
	platform_green_alpha[10][45] = 1'b0; \
	platform_green_alpha[10][46] = 1'b0; \
	platform_green_alpha[10][47] = 1'b0; \
	platform_green_alpha[10][48] = 1'b0; \
	platform_green_alpha[10][49] = 1'b0; \
	platform_green_alpha[10][50] = 1'b0; \
	platform_green_alpha[10][51] = 1'b0; \
	platform_green_alpha[10][52] = 1'b0; \
	platform_green_alpha[10][53] = 1'b0; \
	platform_green_alpha[10][54] = 1'b0; \
	platform_green_alpha[10][55] = 1'b0; \
	platform_green_alpha[10][56] = 1'b0; \
	platform_green_alpha[10][57] = 1'b0; \
	platform_green_alpha[10][58] = 1'b0; \
	platform_green_alpha[10][59] = 1'b0; \
	platform_green_alpha[10][60] = 1'b0; \
	platform_green_alpha[10][61] = 1'b0; \
	platform_green_alpha[10][62] = 1'b0; \
	platform_green_alpha[10][63] = 1'b0; \
	platform_green_alpha[10][64] = 1'b0; \
	platform_green_alpha[10][65] = 1'b0; \
	platform_green_alpha[10][66] = 1'b0; \
	platform_green_alpha[10][67] = 1'b0; \
	platform_green_alpha[10][68] = 1'b0; \
	platform_green_alpha[10][69] = 1'b0; \
	platform_green_alpha[10][70] = 1'b0; \
	platform_green_alpha[10][71] = 1'b0; \
	platform_green_alpha[10][72] = 1'b0; \
	platform_green_alpha[10][73] = 1'b0; \
	platform_green_alpha[10][74] = 1'b0; \
	platform_green_alpha[10][75] = 1'b0; \
	platform_green_alpha[10][76] = 1'b0; \
	platform_green_alpha[10][77] = 1'b0; \
	platform_green_alpha[10][78] = 1'b0; \
	platform_green_alpha[10][79] = 1'b0; \
	platform_green_alpha[10][80] = 1'b0; \
	platform_green_alpha[10][81] = 1'b0; \
	platform_green_alpha[10][82] = 1'b0; \
	platform_green_alpha[10][83] = 1'b0; \
	platform_green_alpha[10][84] = 1'b0; \
	platform_green_alpha[10][85] = 1'b0; \
	platform_green_alpha[10][86] = 1'b0; \
	platform_green_alpha[10][87] = 1'b0; \
	platform_green_alpha[10][88] = 1'b0; \
	platform_green_alpha[10][89] = 1'b0; \
	platform_green_alpha[10][90] = 1'b0; \
	platform_green_alpha[10][91] = 1'b0; \
	platform_green_alpha[10][92] = 1'b0; \
	platform_green_alpha[10][93] = 1'b0; \
	platform_green_alpha[10][94] = 1'b0; \
	platform_green_alpha[10][95] = 1'b1; \
	platform_green_alpha[10][96] = 1'b1; \
	platform_green_alpha[10][97] = 1'b1; \
	platform_green_alpha[10][98] = 1'b1; \
	platform_green_alpha[10][99] = 1'b1; \
	platform_green_alpha[11][0] = 1'b1; \
	platform_green_alpha[11][1] = 1'b1; \
	platform_green_alpha[11][2] = 1'b1; \
	platform_green_alpha[11][3] = 1'b1; \
	platform_green_alpha[11][4] = 1'b1; \
	platform_green_alpha[11][5] = 1'b0; \
	platform_green_alpha[11][6] = 1'b0; \
	platform_green_alpha[11][7] = 1'b0; \
	platform_green_alpha[11][8] = 1'b0; \
	platform_green_alpha[11][9] = 1'b0; \
	platform_green_alpha[11][10] = 1'b0; \
	platform_green_alpha[11][11] = 1'b0; \
	platform_green_alpha[11][12] = 1'b0; \
	platform_green_alpha[11][13] = 1'b0; \
	platform_green_alpha[11][14] = 1'b0; \
	platform_green_alpha[11][15] = 1'b0; \
	platform_green_alpha[11][16] = 1'b0; \
	platform_green_alpha[11][17] = 1'b0; \
	platform_green_alpha[11][18] = 1'b0; \
	platform_green_alpha[11][19] = 1'b0; \
	platform_green_alpha[11][20] = 1'b0; \
	platform_green_alpha[11][21] = 1'b0; \
	platform_green_alpha[11][22] = 1'b0; \
	platform_green_alpha[11][23] = 1'b0; \
	platform_green_alpha[11][24] = 1'b0; \
	platform_green_alpha[11][25] = 1'b0; \
	platform_green_alpha[11][26] = 1'b0; \
	platform_green_alpha[11][27] = 1'b0; \
	platform_green_alpha[11][28] = 1'b0; \
	platform_green_alpha[11][29] = 1'b0; \
	platform_green_alpha[11][30] = 1'b0; \
	platform_green_alpha[11][31] = 1'b0; \
	platform_green_alpha[11][32] = 1'b0; \
	platform_green_alpha[11][33] = 1'b0; \
	platform_green_alpha[11][34] = 1'b0; \
	platform_green_alpha[11][35] = 1'b0; \
	platform_green_alpha[11][36] = 1'b0; \
	platform_green_alpha[11][37] = 1'b0; \
	platform_green_alpha[11][38] = 1'b0; \
	platform_green_alpha[11][39] = 1'b0; \
	platform_green_alpha[11][40] = 1'b0; \
	platform_green_alpha[11][41] = 1'b0; \
	platform_green_alpha[11][42] = 1'b0; \
	platform_green_alpha[11][43] = 1'b0; \
	platform_green_alpha[11][44] = 1'b0; \
	platform_green_alpha[11][45] = 1'b0; \
	platform_green_alpha[11][46] = 1'b0; \
	platform_green_alpha[11][47] = 1'b0; \
	platform_green_alpha[11][48] = 1'b0; \
	platform_green_alpha[11][49] = 1'b0; \
	platform_green_alpha[11][50] = 1'b0; \
	platform_green_alpha[11][51] = 1'b0; \
	platform_green_alpha[11][52] = 1'b0; \
	platform_green_alpha[11][53] = 1'b0; \
	platform_green_alpha[11][54] = 1'b0; \
	platform_green_alpha[11][55] = 1'b0; \
	platform_green_alpha[11][56] = 1'b0; \
	platform_green_alpha[11][57] = 1'b0; \
	platform_green_alpha[11][58] = 1'b0; \
	platform_green_alpha[11][59] = 1'b0; \
	platform_green_alpha[11][60] = 1'b0; \
	platform_green_alpha[11][61] = 1'b0; \
	platform_green_alpha[11][62] = 1'b0; \
	platform_green_alpha[11][63] = 1'b0; \
	platform_green_alpha[11][64] = 1'b0; \
	platform_green_alpha[11][65] = 1'b0; \
	platform_green_alpha[11][66] = 1'b0; \
	platform_green_alpha[11][67] = 1'b0; \
	platform_green_alpha[11][68] = 1'b0; \
	platform_green_alpha[11][69] = 1'b0; \
	platform_green_alpha[11][70] = 1'b0; \
	platform_green_alpha[11][71] = 1'b0; \
	platform_green_alpha[11][72] = 1'b0; \
	platform_green_alpha[11][73] = 1'b0; \
	platform_green_alpha[11][74] = 1'b0; \
	platform_green_alpha[11][75] = 1'b0; \
	platform_green_alpha[11][76] = 1'b0; \
	platform_green_alpha[11][77] = 1'b0; \
	platform_green_alpha[11][78] = 1'b0; \
	platform_green_alpha[11][79] = 1'b0; \
	platform_green_alpha[11][80] = 1'b0; \
	platform_green_alpha[11][81] = 1'b0; \
	platform_green_alpha[11][82] = 1'b0; \
	platform_green_alpha[11][83] = 1'b0; \
	platform_green_alpha[11][84] = 1'b0; \
	platform_green_alpha[11][85] = 1'b0; \
	platform_green_alpha[11][86] = 1'b0; \
	platform_green_alpha[11][87] = 1'b0; \
	platform_green_alpha[11][88] = 1'b0; \
	platform_green_alpha[11][89] = 1'b0; \
	platform_green_alpha[11][90] = 1'b0; \
	platform_green_alpha[11][91] = 1'b0; \
	platform_green_alpha[11][92] = 1'b0; \
	platform_green_alpha[11][93] = 1'b0; \
	platform_green_alpha[11][94] = 1'b0; \
	platform_green_alpha[11][95] = 1'b1; \
	platform_green_alpha[11][96] = 1'b1; \
	platform_green_alpha[11][97] = 1'b1; \
	platform_green_alpha[11][98] = 1'b1; \
	platform_green_alpha[11][99] = 1'b1; \
	platform_green_alpha[12][0] = 1'b1; \
	platform_green_alpha[12][1] = 1'b1; \
	platform_green_alpha[12][2] = 1'b1; \
	platform_green_alpha[12][3] = 1'b1; \
	platform_green_alpha[12][4] = 1'b1; \
	platform_green_alpha[12][5] = 1'b0; \
	platform_green_alpha[12][6] = 1'b0; \
	platform_green_alpha[12][7] = 1'b0; \
	platform_green_alpha[12][8] = 1'b0; \
	platform_green_alpha[12][9] = 1'b0; \
	platform_green_alpha[12][10] = 1'b0; \
	platform_green_alpha[12][11] = 1'b0; \
	platform_green_alpha[12][12] = 1'b0; \
	platform_green_alpha[12][13] = 1'b0; \
	platform_green_alpha[12][14] = 1'b0; \
	platform_green_alpha[12][15] = 1'b0; \
	platform_green_alpha[12][16] = 1'b0; \
	platform_green_alpha[12][17] = 1'b0; \
	platform_green_alpha[12][18] = 1'b0; \
	platform_green_alpha[12][19] = 1'b0; \
	platform_green_alpha[12][20] = 1'b0; \
	platform_green_alpha[12][21] = 1'b0; \
	platform_green_alpha[12][22] = 1'b0; \
	platform_green_alpha[12][23] = 1'b0; \
	platform_green_alpha[12][24] = 1'b0; \
	platform_green_alpha[12][25] = 1'b0; \
	platform_green_alpha[12][26] = 1'b0; \
	platform_green_alpha[12][27] = 1'b0; \
	platform_green_alpha[12][28] = 1'b0; \
	platform_green_alpha[12][29] = 1'b0; \
	platform_green_alpha[12][30] = 1'b0; \
	platform_green_alpha[12][31] = 1'b0; \
	platform_green_alpha[12][32] = 1'b0; \
	platform_green_alpha[12][33] = 1'b0; \
	platform_green_alpha[12][34] = 1'b0; \
	platform_green_alpha[12][35] = 1'b0; \
	platform_green_alpha[12][36] = 1'b0; \
	platform_green_alpha[12][37] = 1'b0; \
	platform_green_alpha[12][38] = 1'b0; \
	platform_green_alpha[12][39] = 1'b0; \
	platform_green_alpha[12][40] = 1'b0; \
	platform_green_alpha[12][41] = 1'b0; \
	platform_green_alpha[12][42] = 1'b0; \
	platform_green_alpha[12][43] = 1'b0; \
	platform_green_alpha[12][44] = 1'b0; \
	platform_green_alpha[12][45] = 1'b0; \
	platform_green_alpha[12][46] = 1'b0; \
	platform_green_alpha[12][47] = 1'b0; \
	platform_green_alpha[12][48] = 1'b0; \
	platform_green_alpha[12][49] = 1'b0; \
	platform_green_alpha[12][50] = 1'b0; \
	platform_green_alpha[12][51] = 1'b0; \
	platform_green_alpha[12][52] = 1'b0; \
	platform_green_alpha[12][53] = 1'b0; \
	platform_green_alpha[12][54] = 1'b0; \
	platform_green_alpha[12][55] = 1'b0; \
	platform_green_alpha[12][56] = 1'b0; \
	platform_green_alpha[12][57] = 1'b0; \
	platform_green_alpha[12][58] = 1'b0; \
	platform_green_alpha[12][59] = 1'b0; \
	platform_green_alpha[12][60] = 1'b0; \
	platform_green_alpha[12][61] = 1'b0; \
	platform_green_alpha[12][62] = 1'b0; \
	platform_green_alpha[12][63] = 1'b0; \
	platform_green_alpha[12][64] = 1'b0; \
	platform_green_alpha[12][65] = 1'b0; \
	platform_green_alpha[12][66] = 1'b0; \
	platform_green_alpha[12][67] = 1'b0; \
	platform_green_alpha[12][68] = 1'b0; \
	platform_green_alpha[12][69] = 1'b0; \
	platform_green_alpha[12][70] = 1'b0; \
	platform_green_alpha[12][71] = 1'b0; \
	platform_green_alpha[12][72] = 1'b0; \
	platform_green_alpha[12][73] = 1'b0; \
	platform_green_alpha[12][74] = 1'b0; \
	platform_green_alpha[12][75] = 1'b0; \
	platform_green_alpha[12][76] = 1'b0; \
	platform_green_alpha[12][77] = 1'b0; \
	platform_green_alpha[12][78] = 1'b0; \
	platform_green_alpha[12][79] = 1'b0; \
	platform_green_alpha[12][80] = 1'b0; \
	platform_green_alpha[12][81] = 1'b0; \
	platform_green_alpha[12][82] = 1'b0; \
	platform_green_alpha[12][83] = 1'b0; \
	platform_green_alpha[12][84] = 1'b0; \
	platform_green_alpha[12][85] = 1'b0; \
	platform_green_alpha[12][86] = 1'b0; \
	platform_green_alpha[12][87] = 1'b0; \
	platform_green_alpha[12][88] = 1'b0; \
	platform_green_alpha[12][89] = 1'b0; \
	platform_green_alpha[12][90] = 1'b0; \
	platform_green_alpha[12][91] = 1'b0; \
	platform_green_alpha[12][92] = 1'b0; \
	platform_green_alpha[12][93] = 1'b0; \
	platform_green_alpha[12][94] = 1'b0; \
	platform_green_alpha[12][95] = 1'b1; \
	platform_green_alpha[12][96] = 1'b1; \
	platform_green_alpha[12][97] = 1'b1; \
	platform_green_alpha[12][98] = 1'b1; \
	platform_green_alpha[12][99] = 1'b1; \
	platform_green_alpha[13][0] = 1'b1; \
	platform_green_alpha[13][1] = 1'b1; \
	platform_green_alpha[13][2] = 1'b1; \
	platform_green_alpha[13][3] = 1'b1; \
	platform_green_alpha[13][4] = 1'b1; \
	platform_green_alpha[13][5] = 1'b0; \
	platform_green_alpha[13][6] = 1'b0; \
	platform_green_alpha[13][7] = 1'b0; \
	platform_green_alpha[13][8] = 1'b0; \
	platform_green_alpha[13][9] = 1'b0; \
	platform_green_alpha[13][10] = 1'b0; \
	platform_green_alpha[13][11] = 1'b0; \
	platform_green_alpha[13][12] = 1'b0; \
	platform_green_alpha[13][13] = 1'b0; \
	platform_green_alpha[13][14] = 1'b0; \
	platform_green_alpha[13][15] = 1'b0; \
	platform_green_alpha[13][16] = 1'b0; \
	platform_green_alpha[13][17] = 1'b0; \
	platform_green_alpha[13][18] = 1'b0; \
	platform_green_alpha[13][19] = 1'b0; \
	platform_green_alpha[13][20] = 1'b0; \
	platform_green_alpha[13][21] = 1'b0; \
	platform_green_alpha[13][22] = 1'b0; \
	platform_green_alpha[13][23] = 1'b0; \
	platform_green_alpha[13][24] = 1'b0; \
	platform_green_alpha[13][25] = 1'b0; \
	platform_green_alpha[13][26] = 1'b0; \
	platform_green_alpha[13][27] = 1'b0; \
	platform_green_alpha[13][28] = 1'b0; \
	platform_green_alpha[13][29] = 1'b0; \
	platform_green_alpha[13][30] = 1'b0; \
	platform_green_alpha[13][31] = 1'b0; \
	platform_green_alpha[13][32] = 1'b0; \
	platform_green_alpha[13][33] = 1'b0; \
	platform_green_alpha[13][34] = 1'b0; \
	platform_green_alpha[13][35] = 1'b0; \
	platform_green_alpha[13][36] = 1'b0; \
	platform_green_alpha[13][37] = 1'b0; \
	platform_green_alpha[13][38] = 1'b0; \
	platform_green_alpha[13][39] = 1'b0; \
	platform_green_alpha[13][40] = 1'b0; \
	platform_green_alpha[13][41] = 1'b0; \
	platform_green_alpha[13][42] = 1'b0; \
	platform_green_alpha[13][43] = 1'b0; \
	platform_green_alpha[13][44] = 1'b0; \
	platform_green_alpha[13][45] = 1'b0; \
	platform_green_alpha[13][46] = 1'b0; \
	platform_green_alpha[13][47] = 1'b0; \
	platform_green_alpha[13][48] = 1'b0; \
	platform_green_alpha[13][49] = 1'b0; \
	platform_green_alpha[13][50] = 1'b0; \
	platform_green_alpha[13][51] = 1'b0; \
	platform_green_alpha[13][52] = 1'b0; \
	platform_green_alpha[13][53] = 1'b0; \
	platform_green_alpha[13][54] = 1'b0; \
	platform_green_alpha[13][55] = 1'b0; \
	platform_green_alpha[13][56] = 1'b0; \
	platform_green_alpha[13][57] = 1'b0; \
	platform_green_alpha[13][58] = 1'b0; \
	platform_green_alpha[13][59] = 1'b0; \
	platform_green_alpha[13][60] = 1'b0; \
	platform_green_alpha[13][61] = 1'b0; \
	platform_green_alpha[13][62] = 1'b0; \
	platform_green_alpha[13][63] = 1'b0; \
	platform_green_alpha[13][64] = 1'b0; \
	platform_green_alpha[13][65] = 1'b0; \
	platform_green_alpha[13][66] = 1'b0; \
	platform_green_alpha[13][67] = 1'b0; \
	platform_green_alpha[13][68] = 1'b0; \
	platform_green_alpha[13][69] = 1'b0; \
	platform_green_alpha[13][70] = 1'b0; \
	platform_green_alpha[13][71] = 1'b0; \
	platform_green_alpha[13][72] = 1'b0; \
	platform_green_alpha[13][73] = 1'b0; \
	platform_green_alpha[13][74] = 1'b0; \
	platform_green_alpha[13][75] = 1'b0; \
	platform_green_alpha[13][76] = 1'b0; \
	platform_green_alpha[13][77] = 1'b0; \
	platform_green_alpha[13][78] = 1'b0; \
	platform_green_alpha[13][79] = 1'b0; \
	platform_green_alpha[13][80] = 1'b0; \
	platform_green_alpha[13][81] = 1'b0; \
	platform_green_alpha[13][82] = 1'b0; \
	platform_green_alpha[13][83] = 1'b0; \
	platform_green_alpha[13][84] = 1'b0; \
	platform_green_alpha[13][85] = 1'b0; \
	platform_green_alpha[13][86] = 1'b0; \
	platform_green_alpha[13][87] = 1'b0; \
	platform_green_alpha[13][88] = 1'b0; \
	platform_green_alpha[13][89] = 1'b0; \
	platform_green_alpha[13][90] = 1'b0; \
	platform_green_alpha[13][91] = 1'b0; \
	platform_green_alpha[13][92] = 1'b0; \
	platform_green_alpha[13][93] = 1'b0; \
	platform_green_alpha[13][94] = 1'b0; \
	platform_green_alpha[13][95] = 1'b1; \
	platform_green_alpha[13][96] = 1'b1; \
	platform_green_alpha[13][97] = 1'b1; \
	platform_green_alpha[13][98] = 1'b1; \
	platform_green_alpha[13][99] = 1'b1; \
	platform_green_alpha[14][0] = 1'b1; \
	platform_green_alpha[14][1] = 1'b1; \
	platform_green_alpha[14][2] = 1'b1; \
	platform_green_alpha[14][3] = 1'b1; \
	platform_green_alpha[14][4] = 1'b1; \
	platform_green_alpha[14][5] = 1'b0; \
	platform_green_alpha[14][6] = 1'b0; \
	platform_green_alpha[14][7] = 1'b0; \
	platform_green_alpha[14][8] = 1'b0; \
	platform_green_alpha[14][9] = 1'b0; \
	platform_green_alpha[14][10] = 1'b0; \
	platform_green_alpha[14][11] = 1'b0; \
	platform_green_alpha[14][12] = 1'b0; \
	platform_green_alpha[14][13] = 1'b0; \
	platform_green_alpha[14][14] = 1'b0; \
	platform_green_alpha[14][15] = 1'b0; \
	platform_green_alpha[14][16] = 1'b0; \
	platform_green_alpha[14][17] = 1'b0; \
	platform_green_alpha[14][18] = 1'b0; \
	platform_green_alpha[14][19] = 1'b0; \
	platform_green_alpha[14][20] = 1'b0; \
	platform_green_alpha[14][21] = 1'b0; \
	platform_green_alpha[14][22] = 1'b0; \
	platform_green_alpha[14][23] = 1'b0; \
	platform_green_alpha[14][24] = 1'b0; \
	platform_green_alpha[14][25] = 1'b0; \
	platform_green_alpha[14][26] = 1'b0; \
	platform_green_alpha[14][27] = 1'b0; \
	platform_green_alpha[14][28] = 1'b0; \
	platform_green_alpha[14][29] = 1'b0; \
	platform_green_alpha[14][30] = 1'b0; \
	platform_green_alpha[14][31] = 1'b0; \
	platform_green_alpha[14][32] = 1'b0; \
	platform_green_alpha[14][33] = 1'b0; \
	platform_green_alpha[14][34] = 1'b0; \
	platform_green_alpha[14][35] = 1'b0; \
	platform_green_alpha[14][36] = 1'b0; \
	platform_green_alpha[14][37] = 1'b0; \
	platform_green_alpha[14][38] = 1'b0; \
	platform_green_alpha[14][39] = 1'b0; \
	platform_green_alpha[14][40] = 1'b0; \
	platform_green_alpha[14][41] = 1'b0; \
	platform_green_alpha[14][42] = 1'b0; \
	platform_green_alpha[14][43] = 1'b0; \
	platform_green_alpha[14][44] = 1'b0; \
	platform_green_alpha[14][45] = 1'b0; \
	platform_green_alpha[14][46] = 1'b0; \
	platform_green_alpha[14][47] = 1'b0; \
	platform_green_alpha[14][48] = 1'b0; \
	platform_green_alpha[14][49] = 1'b0; \
	platform_green_alpha[14][50] = 1'b0; \
	platform_green_alpha[14][51] = 1'b0; \
	platform_green_alpha[14][52] = 1'b0; \
	platform_green_alpha[14][53] = 1'b0; \
	platform_green_alpha[14][54] = 1'b0; \
	platform_green_alpha[14][55] = 1'b0; \
	platform_green_alpha[14][56] = 1'b0; \
	platform_green_alpha[14][57] = 1'b0; \
	platform_green_alpha[14][58] = 1'b0; \
	platform_green_alpha[14][59] = 1'b0; \
	platform_green_alpha[14][60] = 1'b0; \
	platform_green_alpha[14][61] = 1'b0; \
	platform_green_alpha[14][62] = 1'b0; \
	platform_green_alpha[14][63] = 1'b0; \
	platform_green_alpha[14][64] = 1'b0; \
	platform_green_alpha[14][65] = 1'b0; \
	platform_green_alpha[14][66] = 1'b0; \
	platform_green_alpha[14][67] = 1'b0; \
	platform_green_alpha[14][68] = 1'b0; \
	platform_green_alpha[14][69] = 1'b0; \
	platform_green_alpha[14][70] = 1'b0; \
	platform_green_alpha[14][71] = 1'b0; \
	platform_green_alpha[14][72] = 1'b0; \
	platform_green_alpha[14][73] = 1'b0; \
	platform_green_alpha[14][74] = 1'b0; \
	platform_green_alpha[14][75] = 1'b0; \
	platform_green_alpha[14][76] = 1'b0; \
	platform_green_alpha[14][77] = 1'b0; \
	platform_green_alpha[14][78] = 1'b0; \
	platform_green_alpha[14][79] = 1'b0; \
	platform_green_alpha[14][80] = 1'b0; \
	platform_green_alpha[14][81] = 1'b0; \
	platform_green_alpha[14][82] = 1'b0; \
	platform_green_alpha[14][83] = 1'b0; \
	platform_green_alpha[14][84] = 1'b0; \
	platform_green_alpha[14][85] = 1'b0; \
	platform_green_alpha[14][86] = 1'b0; \
	platform_green_alpha[14][87] = 1'b0; \
	platform_green_alpha[14][88] = 1'b0; \
	platform_green_alpha[14][89] = 1'b0; \
	platform_green_alpha[14][90] = 1'b0; \
	platform_green_alpha[14][91] = 1'b0; \
	platform_green_alpha[14][92] = 1'b0; \
	platform_green_alpha[14][93] = 1'b0; \
	platform_green_alpha[14][94] = 1'b0; \
	platform_green_alpha[14][95] = 1'b1; \
	platform_green_alpha[14][96] = 1'b1; \
	platform_green_alpha[14][97] = 1'b1; \
	platform_green_alpha[14][98] = 1'b1; \
	platform_green_alpha[14][99] = 1'b1; \
	platform_green_alpha[15][0] = 1'b1; \
	platform_green_alpha[15][1] = 1'b1; \
	platform_green_alpha[15][2] = 1'b1; \
	platform_green_alpha[15][3] = 1'b1; \
	platform_green_alpha[15][4] = 1'b1; \
	platform_green_alpha[15][5] = 1'b0; \
	platform_green_alpha[15][6] = 1'b0; \
	platform_green_alpha[15][7] = 1'b0; \
	platform_green_alpha[15][8] = 1'b0; \
	platform_green_alpha[15][9] = 1'b0; \
	platform_green_alpha[15][10] = 1'b0; \
	platform_green_alpha[15][11] = 1'b0; \
	platform_green_alpha[15][12] = 1'b0; \
	platform_green_alpha[15][13] = 1'b0; \
	platform_green_alpha[15][14] = 1'b0; \
	platform_green_alpha[15][15] = 1'b0; \
	platform_green_alpha[15][16] = 1'b0; \
	platform_green_alpha[15][17] = 1'b0; \
	platform_green_alpha[15][18] = 1'b0; \
	platform_green_alpha[15][19] = 1'b0; \
	platform_green_alpha[15][20] = 1'b0; \
	platform_green_alpha[15][21] = 1'b0; \
	platform_green_alpha[15][22] = 1'b0; \
	platform_green_alpha[15][23] = 1'b0; \
	platform_green_alpha[15][24] = 1'b0; \
	platform_green_alpha[15][25] = 1'b0; \
	platform_green_alpha[15][26] = 1'b0; \
	platform_green_alpha[15][27] = 1'b0; \
	platform_green_alpha[15][28] = 1'b0; \
	platform_green_alpha[15][29] = 1'b0; \
	platform_green_alpha[15][30] = 1'b0; \
	platform_green_alpha[15][31] = 1'b0; \
	platform_green_alpha[15][32] = 1'b0; \
	platform_green_alpha[15][33] = 1'b0; \
	platform_green_alpha[15][34] = 1'b0; \
	platform_green_alpha[15][35] = 1'b0; \
	platform_green_alpha[15][36] = 1'b0; \
	platform_green_alpha[15][37] = 1'b0; \
	platform_green_alpha[15][38] = 1'b0; \
	platform_green_alpha[15][39] = 1'b0; \
	platform_green_alpha[15][40] = 1'b0; \
	platform_green_alpha[15][41] = 1'b0; \
	platform_green_alpha[15][42] = 1'b0; \
	platform_green_alpha[15][43] = 1'b0; \
	platform_green_alpha[15][44] = 1'b0; \
	platform_green_alpha[15][45] = 1'b0; \
	platform_green_alpha[15][46] = 1'b0; \
	platform_green_alpha[15][47] = 1'b0; \
	platform_green_alpha[15][48] = 1'b0; \
	platform_green_alpha[15][49] = 1'b0; \
	platform_green_alpha[15][50] = 1'b0; \
	platform_green_alpha[15][51] = 1'b0; \
	platform_green_alpha[15][52] = 1'b0; \
	platform_green_alpha[15][53] = 1'b0; \
	platform_green_alpha[15][54] = 1'b0; \
	platform_green_alpha[15][55] = 1'b0; \
	platform_green_alpha[15][56] = 1'b0; \
	platform_green_alpha[15][57] = 1'b0; \
	platform_green_alpha[15][58] = 1'b0; \
	platform_green_alpha[15][59] = 1'b0; \
	platform_green_alpha[15][60] = 1'b0; \
	platform_green_alpha[15][61] = 1'b0; \
	platform_green_alpha[15][62] = 1'b0; \
	platform_green_alpha[15][63] = 1'b0; \
	platform_green_alpha[15][64] = 1'b0; \
	platform_green_alpha[15][65] = 1'b0; \
	platform_green_alpha[15][66] = 1'b0; \
	platform_green_alpha[15][67] = 1'b0; \
	platform_green_alpha[15][68] = 1'b0; \
	platform_green_alpha[15][69] = 1'b0; \
	platform_green_alpha[15][70] = 1'b0; \
	platform_green_alpha[15][71] = 1'b0; \
	platform_green_alpha[15][72] = 1'b0; \
	platform_green_alpha[15][73] = 1'b0; \
	platform_green_alpha[15][74] = 1'b0; \
	platform_green_alpha[15][75] = 1'b0; \
	platform_green_alpha[15][76] = 1'b0; \
	platform_green_alpha[15][77] = 1'b0; \
	platform_green_alpha[15][78] = 1'b0; \
	platform_green_alpha[15][79] = 1'b0; \
	platform_green_alpha[15][80] = 1'b0; \
	platform_green_alpha[15][81] = 1'b0; \
	platform_green_alpha[15][82] = 1'b0; \
	platform_green_alpha[15][83] = 1'b0; \
	platform_green_alpha[15][84] = 1'b0; \
	platform_green_alpha[15][85] = 1'b0; \
	platform_green_alpha[15][86] = 1'b0; \
	platform_green_alpha[15][87] = 1'b0; \
	platform_green_alpha[15][88] = 1'b0; \
	platform_green_alpha[15][89] = 1'b0; \
	platform_green_alpha[15][90] = 1'b0; \
	platform_green_alpha[15][91] = 1'b0; \
	platform_green_alpha[15][92] = 1'b0; \
	platform_green_alpha[15][93] = 1'b0; \
	platform_green_alpha[15][94] = 1'b0; \
	platform_green_alpha[15][95] = 1'b1; \
	platform_green_alpha[15][96] = 1'b1; \
	platform_green_alpha[15][97] = 1'b1; \
	platform_green_alpha[15][98] = 1'b1; \
	platform_green_alpha[15][99] = 1'b1; \
	platform_green_alpha[16][0] = 1'b1; \
	platform_green_alpha[16][1] = 1'b1; \
	platform_green_alpha[16][2] = 1'b1; \
	platform_green_alpha[16][3] = 1'b1; \
	platform_green_alpha[16][4] = 1'b1; \
	platform_green_alpha[16][5] = 1'b0; \
	platform_green_alpha[16][6] = 1'b0; \
	platform_green_alpha[16][7] = 1'b0; \
	platform_green_alpha[16][8] = 1'b0; \
	platform_green_alpha[16][9] = 1'b0; \
	platform_green_alpha[16][10] = 1'b0; \
	platform_green_alpha[16][11] = 1'b0; \
	platform_green_alpha[16][12] = 1'b0; \
	platform_green_alpha[16][13] = 1'b0; \
	platform_green_alpha[16][14] = 1'b0; \
	platform_green_alpha[16][15] = 1'b0; \
	platform_green_alpha[16][16] = 1'b0; \
	platform_green_alpha[16][17] = 1'b0; \
	platform_green_alpha[16][18] = 1'b0; \
	platform_green_alpha[16][19] = 1'b0; \
	platform_green_alpha[16][20] = 1'b0; \
	platform_green_alpha[16][21] = 1'b0; \
	platform_green_alpha[16][22] = 1'b0; \
	platform_green_alpha[16][23] = 1'b0; \
	platform_green_alpha[16][24] = 1'b0; \
	platform_green_alpha[16][25] = 1'b0; \
	platform_green_alpha[16][26] = 1'b0; \
	platform_green_alpha[16][27] = 1'b0; \
	platform_green_alpha[16][28] = 1'b0; \
	platform_green_alpha[16][29] = 1'b0; \
	platform_green_alpha[16][30] = 1'b0; \
	platform_green_alpha[16][31] = 1'b0; \
	platform_green_alpha[16][32] = 1'b0; \
	platform_green_alpha[16][33] = 1'b0; \
	platform_green_alpha[16][34] = 1'b0; \
	platform_green_alpha[16][35] = 1'b0; \
	platform_green_alpha[16][36] = 1'b0; \
	platform_green_alpha[16][37] = 1'b0; \
	platform_green_alpha[16][38] = 1'b0; \
	platform_green_alpha[16][39] = 1'b0; \
	platform_green_alpha[16][40] = 1'b0; \
	platform_green_alpha[16][41] = 1'b0; \
	platform_green_alpha[16][42] = 1'b0; \
	platform_green_alpha[16][43] = 1'b0; \
	platform_green_alpha[16][44] = 1'b0; \
	platform_green_alpha[16][45] = 1'b0; \
	platform_green_alpha[16][46] = 1'b0; \
	platform_green_alpha[16][47] = 1'b0; \
	platform_green_alpha[16][48] = 1'b0; \
	platform_green_alpha[16][49] = 1'b0; \
	platform_green_alpha[16][50] = 1'b0; \
	platform_green_alpha[16][51] = 1'b0; \
	platform_green_alpha[16][52] = 1'b0; \
	platform_green_alpha[16][53] = 1'b0; \
	platform_green_alpha[16][54] = 1'b0; \
	platform_green_alpha[16][55] = 1'b0; \
	platform_green_alpha[16][56] = 1'b0; \
	platform_green_alpha[16][57] = 1'b0; \
	platform_green_alpha[16][58] = 1'b0; \
	platform_green_alpha[16][59] = 1'b0; \
	platform_green_alpha[16][60] = 1'b0; \
	platform_green_alpha[16][61] = 1'b0; \
	platform_green_alpha[16][62] = 1'b0; \
	platform_green_alpha[16][63] = 1'b0; \
	platform_green_alpha[16][64] = 1'b0; \
	platform_green_alpha[16][65] = 1'b0; \
	platform_green_alpha[16][66] = 1'b0; \
	platform_green_alpha[16][67] = 1'b0; \
	platform_green_alpha[16][68] = 1'b0; \
	platform_green_alpha[16][69] = 1'b0; \
	platform_green_alpha[16][70] = 1'b0; \
	platform_green_alpha[16][71] = 1'b0; \
	platform_green_alpha[16][72] = 1'b0; \
	platform_green_alpha[16][73] = 1'b0; \
	platform_green_alpha[16][74] = 1'b0; \
	platform_green_alpha[16][75] = 1'b0; \
	platform_green_alpha[16][76] = 1'b0; \
	platform_green_alpha[16][77] = 1'b0; \
	platform_green_alpha[16][78] = 1'b0; \
	platform_green_alpha[16][79] = 1'b0; \
	platform_green_alpha[16][80] = 1'b0; \
	platform_green_alpha[16][81] = 1'b0; \
	platform_green_alpha[16][82] = 1'b0; \
	platform_green_alpha[16][83] = 1'b0; \
	platform_green_alpha[16][84] = 1'b0; \
	platform_green_alpha[16][85] = 1'b0; \
	platform_green_alpha[16][86] = 1'b0; \
	platform_green_alpha[16][87] = 1'b0; \
	platform_green_alpha[16][88] = 1'b0; \
	platform_green_alpha[16][89] = 1'b0; \
	platform_green_alpha[16][90] = 1'b0; \
	platform_green_alpha[16][91] = 1'b0; \
	platform_green_alpha[16][92] = 1'b0; \
	platform_green_alpha[16][93] = 1'b0; \
	platform_green_alpha[16][94] = 1'b0; \
	platform_green_alpha[16][95] = 1'b1; \
	platform_green_alpha[16][96] = 1'b1; \
	platform_green_alpha[16][97] = 1'b1; \
	platform_green_alpha[16][98] = 1'b1; \
	platform_green_alpha[16][99] = 1'b1; \
	platform_green_alpha[17][0] = 1'b1; \
	platform_green_alpha[17][1] = 1'b1; \
	platform_green_alpha[17][2] = 1'b1; \
	platform_green_alpha[17][3] = 1'b1; \
	platform_green_alpha[17][4] = 1'b1; \
	platform_green_alpha[17][5] = 1'b0; \
	platform_green_alpha[17][6] = 1'b0; \
	platform_green_alpha[17][7] = 1'b0; \
	platform_green_alpha[17][8] = 1'b0; \
	platform_green_alpha[17][9] = 1'b0; \
	platform_green_alpha[17][10] = 1'b0; \
	platform_green_alpha[17][11] = 1'b0; \
	platform_green_alpha[17][12] = 1'b0; \
	platform_green_alpha[17][13] = 1'b0; \
	platform_green_alpha[17][14] = 1'b0; \
	platform_green_alpha[17][15] = 1'b0; \
	platform_green_alpha[17][16] = 1'b0; \
	platform_green_alpha[17][17] = 1'b0; \
	platform_green_alpha[17][18] = 1'b0; \
	platform_green_alpha[17][19] = 1'b0; \
	platform_green_alpha[17][20] = 1'b0; \
	platform_green_alpha[17][21] = 1'b0; \
	platform_green_alpha[17][22] = 1'b0; \
	platform_green_alpha[17][23] = 1'b0; \
	platform_green_alpha[17][24] = 1'b0; \
	platform_green_alpha[17][25] = 1'b0; \
	platform_green_alpha[17][26] = 1'b0; \
	platform_green_alpha[17][27] = 1'b0; \
	platform_green_alpha[17][28] = 1'b0; \
	platform_green_alpha[17][29] = 1'b0; \
	platform_green_alpha[17][30] = 1'b0; \
	platform_green_alpha[17][31] = 1'b0; \
	platform_green_alpha[17][32] = 1'b0; \
	platform_green_alpha[17][33] = 1'b0; \
	platform_green_alpha[17][34] = 1'b0; \
	platform_green_alpha[17][35] = 1'b0; \
	platform_green_alpha[17][36] = 1'b0; \
	platform_green_alpha[17][37] = 1'b0; \
	platform_green_alpha[17][38] = 1'b0; \
	platform_green_alpha[17][39] = 1'b0; \
	platform_green_alpha[17][40] = 1'b0; \
	platform_green_alpha[17][41] = 1'b0; \
	platform_green_alpha[17][42] = 1'b0; \
	platform_green_alpha[17][43] = 1'b0; \
	platform_green_alpha[17][44] = 1'b0; \
	platform_green_alpha[17][45] = 1'b0; \
	platform_green_alpha[17][46] = 1'b0; \
	platform_green_alpha[17][47] = 1'b0; \
	platform_green_alpha[17][48] = 1'b0; \
	platform_green_alpha[17][49] = 1'b0; \
	platform_green_alpha[17][50] = 1'b0; \
	platform_green_alpha[17][51] = 1'b0; \
	platform_green_alpha[17][52] = 1'b0; \
	platform_green_alpha[17][53] = 1'b0; \
	platform_green_alpha[17][54] = 1'b0; \
	platform_green_alpha[17][55] = 1'b0; \
	platform_green_alpha[17][56] = 1'b0; \
	platform_green_alpha[17][57] = 1'b0; \
	platform_green_alpha[17][58] = 1'b0; \
	platform_green_alpha[17][59] = 1'b0; \
	platform_green_alpha[17][60] = 1'b0; \
	platform_green_alpha[17][61] = 1'b0; \
	platform_green_alpha[17][62] = 1'b0; \
	platform_green_alpha[17][63] = 1'b0; \
	platform_green_alpha[17][64] = 1'b0; \
	platform_green_alpha[17][65] = 1'b0; \
	platform_green_alpha[17][66] = 1'b0; \
	platform_green_alpha[17][67] = 1'b0; \
	platform_green_alpha[17][68] = 1'b0; \
	platform_green_alpha[17][69] = 1'b0; \
	platform_green_alpha[17][70] = 1'b0; \
	platform_green_alpha[17][71] = 1'b0; \
	platform_green_alpha[17][72] = 1'b0; \
	platform_green_alpha[17][73] = 1'b0; \
	platform_green_alpha[17][74] = 1'b0; \
	platform_green_alpha[17][75] = 1'b0; \
	platform_green_alpha[17][76] = 1'b0; \
	platform_green_alpha[17][77] = 1'b0; \
	platform_green_alpha[17][78] = 1'b0; \
	platform_green_alpha[17][79] = 1'b0; \
	platform_green_alpha[17][80] = 1'b0; \
	platform_green_alpha[17][81] = 1'b0; \
	platform_green_alpha[17][82] = 1'b0; \
	platform_green_alpha[17][83] = 1'b0; \
	platform_green_alpha[17][84] = 1'b0; \
	platform_green_alpha[17][85] = 1'b0; \
	platform_green_alpha[17][86] = 1'b0; \
	platform_green_alpha[17][87] = 1'b0; \
	platform_green_alpha[17][88] = 1'b0; \
	platform_green_alpha[17][89] = 1'b0; \
	platform_green_alpha[17][90] = 1'b0; \
	platform_green_alpha[17][91] = 1'b0; \
	platform_green_alpha[17][92] = 1'b0; \
	platform_green_alpha[17][93] = 1'b0; \
	platform_green_alpha[17][94] = 1'b0; \
	platform_green_alpha[17][95] = 1'b1; \
	platform_green_alpha[17][96] = 1'b1; \
	platform_green_alpha[17][97] = 1'b1; \
	platform_green_alpha[17][98] = 1'b1; \
	platform_green_alpha[17][99] = 1'b1; \
	platform_green_alpha[18][0] = 1'b1; \
	platform_green_alpha[18][1] = 1'b1; \
	platform_green_alpha[18][2] = 1'b1; \
	platform_green_alpha[18][3] = 1'b1; \
	platform_green_alpha[18][4] = 1'b1; \
	platform_green_alpha[18][5] = 1'b0; \
	platform_green_alpha[18][6] = 1'b0; \
	platform_green_alpha[18][7] = 1'b0; \
	platform_green_alpha[18][8] = 1'b0; \
	platform_green_alpha[18][9] = 1'b0; \
	platform_green_alpha[18][10] = 1'b0; \
	platform_green_alpha[18][11] = 1'b0; \
	platform_green_alpha[18][12] = 1'b0; \
	platform_green_alpha[18][13] = 1'b0; \
	platform_green_alpha[18][14] = 1'b0; \
	platform_green_alpha[18][15] = 1'b0; \
	platform_green_alpha[18][16] = 1'b0; \
	platform_green_alpha[18][17] = 1'b0; \
	platform_green_alpha[18][18] = 1'b0; \
	platform_green_alpha[18][19] = 1'b0; \
	platform_green_alpha[18][20] = 1'b0; \
	platform_green_alpha[18][21] = 1'b0; \
	platform_green_alpha[18][22] = 1'b0; \
	platform_green_alpha[18][23] = 1'b0; \
	platform_green_alpha[18][24] = 1'b0; \
	platform_green_alpha[18][25] = 1'b0; \
	platform_green_alpha[18][26] = 1'b0; \
	platform_green_alpha[18][27] = 1'b0; \
	platform_green_alpha[18][28] = 1'b0; \
	platform_green_alpha[18][29] = 1'b0; \
	platform_green_alpha[18][30] = 1'b0; \
	platform_green_alpha[18][31] = 1'b0; \
	platform_green_alpha[18][32] = 1'b0; \
	platform_green_alpha[18][33] = 1'b0; \
	platform_green_alpha[18][34] = 1'b0; \
	platform_green_alpha[18][35] = 1'b0; \
	platform_green_alpha[18][36] = 1'b0; \
	platform_green_alpha[18][37] = 1'b0; \
	platform_green_alpha[18][38] = 1'b0; \
	platform_green_alpha[18][39] = 1'b0; \
	platform_green_alpha[18][40] = 1'b0; \
	platform_green_alpha[18][41] = 1'b0; \
	platform_green_alpha[18][42] = 1'b0; \
	platform_green_alpha[18][43] = 1'b0; \
	platform_green_alpha[18][44] = 1'b0; \
	platform_green_alpha[18][45] = 1'b0; \
	platform_green_alpha[18][46] = 1'b0; \
	platform_green_alpha[18][47] = 1'b0; \
	platform_green_alpha[18][48] = 1'b0; \
	platform_green_alpha[18][49] = 1'b0; \
	platform_green_alpha[18][50] = 1'b0; \
	platform_green_alpha[18][51] = 1'b0; \
	platform_green_alpha[18][52] = 1'b0; \
	platform_green_alpha[18][53] = 1'b0; \
	platform_green_alpha[18][54] = 1'b0; \
	platform_green_alpha[18][55] = 1'b0; \
	platform_green_alpha[18][56] = 1'b0; \
	platform_green_alpha[18][57] = 1'b0; \
	platform_green_alpha[18][58] = 1'b0; \
	platform_green_alpha[18][59] = 1'b0; \
	platform_green_alpha[18][60] = 1'b0; \
	platform_green_alpha[18][61] = 1'b0; \
	platform_green_alpha[18][62] = 1'b0; \
	platform_green_alpha[18][63] = 1'b0; \
	platform_green_alpha[18][64] = 1'b0; \
	platform_green_alpha[18][65] = 1'b0; \
	platform_green_alpha[18][66] = 1'b0; \
	platform_green_alpha[18][67] = 1'b0; \
	platform_green_alpha[18][68] = 1'b0; \
	platform_green_alpha[18][69] = 1'b0; \
	platform_green_alpha[18][70] = 1'b0; \
	platform_green_alpha[18][71] = 1'b0; \
	platform_green_alpha[18][72] = 1'b0; \
	platform_green_alpha[18][73] = 1'b0; \
	platform_green_alpha[18][74] = 1'b0; \
	platform_green_alpha[18][75] = 1'b0; \
	platform_green_alpha[18][76] = 1'b0; \
	platform_green_alpha[18][77] = 1'b0; \
	platform_green_alpha[18][78] = 1'b0; \
	platform_green_alpha[18][79] = 1'b0; \
	platform_green_alpha[18][80] = 1'b0; \
	platform_green_alpha[18][81] = 1'b0; \
	platform_green_alpha[18][82] = 1'b0; \
	platform_green_alpha[18][83] = 1'b0; \
	platform_green_alpha[18][84] = 1'b0; \
	platform_green_alpha[18][85] = 1'b0; \
	platform_green_alpha[18][86] = 1'b0; \
	platform_green_alpha[18][87] = 1'b0; \
	platform_green_alpha[18][88] = 1'b0; \
	platform_green_alpha[18][89] = 1'b0; \
	platform_green_alpha[18][90] = 1'b0; \
	platform_green_alpha[18][91] = 1'b0; \
	platform_green_alpha[18][92] = 1'b0; \
	platform_green_alpha[18][93] = 1'b0; \
	platform_green_alpha[18][94] = 1'b0; \
	platform_green_alpha[18][95] = 1'b1; \
	platform_green_alpha[18][96] = 1'b1; \
	platform_green_alpha[18][97] = 1'b1; \
	platform_green_alpha[18][98] = 1'b1; \
	platform_green_alpha[18][99] = 1'b1; \
	platform_green_alpha[19][0] = 1'b1; \
	platform_green_alpha[19][1] = 1'b1; \
	platform_green_alpha[19][2] = 1'b1; \
	platform_green_alpha[19][3] = 1'b1; \
	platform_green_alpha[19][4] = 1'b1; \
	platform_green_alpha[19][5] = 1'b0; \
	platform_green_alpha[19][6] = 1'b0; \
	platform_green_alpha[19][7] = 1'b0; \
	platform_green_alpha[19][8] = 1'b0; \
	platform_green_alpha[19][9] = 1'b0; \
	platform_green_alpha[19][10] = 1'b0; \
	platform_green_alpha[19][11] = 1'b0; \
	platform_green_alpha[19][12] = 1'b0; \
	platform_green_alpha[19][13] = 1'b0; \
	platform_green_alpha[19][14] = 1'b0; \
	platform_green_alpha[19][15] = 1'b0; \
	platform_green_alpha[19][16] = 1'b0; \
	platform_green_alpha[19][17] = 1'b0; \
	platform_green_alpha[19][18] = 1'b0; \
	platform_green_alpha[19][19] = 1'b0; \
	platform_green_alpha[19][20] = 1'b0; \
	platform_green_alpha[19][21] = 1'b0; \
	platform_green_alpha[19][22] = 1'b0; \
	platform_green_alpha[19][23] = 1'b0; \
	platform_green_alpha[19][24] = 1'b0; \
	platform_green_alpha[19][25] = 1'b0; \
	platform_green_alpha[19][26] = 1'b0; \
	platform_green_alpha[19][27] = 1'b0; \
	platform_green_alpha[19][28] = 1'b0; \
	platform_green_alpha[19][29] = 1'b0; \
	platform_green_alpha[19][30] = 1'b0; \
	platform_green_alpha[19][31] = 1'b0; \
	platform_green_alpha[19][32] = 1'b0; \
	platform_green_alpha[19][33] = 1'b0; \
	platform_green_alpha[19][34] = 1'b0; \
	platform_green_alpha[19][35] = 1'b0; \
	platform_green_alpha[19][36] = 1'b0; \
	platform_green_alpha[19][37] = 1'b0; \
	platform_green_alpha[19][38] = 1'b0; \
	platform_green_alpha[19][39] = 1'b0; \
	platform_green_alpha[19][40] = 1'b0; \
	platform_green_alpha[19][41] = 1'b0; \
	platform_green_alpha[19][42] = 1'b0; \
	platform_green_alpha[19][43] = 1'b0; \
	platform_green_alpha[19][44] = 1'b0; \
	platform_green_alpha[19][45] = 1'b0; \
	platform_green_alpha[19][46] = 1'b0; \
	platform_green_alpha[19][47] = 1'b0; \
	platform_green_alpha[19][48] = 1'b0; \
	platform_green_alpha[19][49] = 1'b0; \
	platform_green_alpha[19][50] = 1'b0; \
	platform_green_alpha[19][51] = 1'b0; \
	platform_green_alpha[19][52] = 1'b0; \
	platform_green_alpha[19][53] = 1'b0; \
	platform_green_alpha[19][54] = 1'b0; \
	platform_green_alpha[19][55] = 1'b0; \
	platform_green_alpha[19][56] = 1'b0; \
	platform_green_alpha[19][57] = 1'b0; \
	platform_green_alpha[19][58] = 1'b0; \
	platform_green_alpha[19][59] = 1'b0; \
	platform_green_alpha[19][60] = 1'b0; \
	platform_green_alpha[19][61] = 1'b0; \
	platform_green_alpha[19][62] = 1'b0; \
	platform_green_alpha[19][63] = 1'b0; \
	platform_green_alpha[19][64] = 1'b0; \
	platform_green_alpha[19][65] = 1'b0; \
	platform_green_alpha[19][66] = 1'b0; \
	platform_green_alpha[19][67] = 1'b0; \
	platform_green_alpha[19][68] = 1'b0; \
	platform_green_alpha[19][69] = 1'b0; \
	platform_green_alpha[19][70] = 1'b0; \
	platform_green_alpha[19][71] = 1'b0; \
	platform_green_alpha[19][72] = 1'b0; \
	platform_green_alpha[19][73] = 1'b0; \
	platform_green_alpha[19][74] = 1'b0; \
	platform_green_alpha[19][75] = 1'b0; \
	platform_green_alpha[19][76] = 1'b0; \
	platform_green_alpha[19][77] = 1'b0; \
	platform_green_alpha[19][78] = 1'b0; \
	platform_green_alpha[19][79] = 1'b0; \
	platform_green_alpha[19][80] = 1'b0; \
	platform_green_alpha[19][81] = 1'b0; \
	platform_green_alpha[19][82] = 1'b0; \
	platform_green_alpha[19][83] = 1'b0; \
	platform_green_alpha[19][84] = 1'b0; \
	platform_green_alpha[19][85] = 1'b0; \
	platform_green_alpha[19][86] = 1'b0; \
	platform_green_alpha[19][87] = 1'b0; \
	platform_green_alpha[19][88] = 1'b0; \
	platform_green_alpha[19][89] = 1'b0; \
	platform_green_alpha[19][90] = 1'b0; \
	platform_green_alpha[19][91] = 1'b0; \
	platform_green_alpha[19][92] = 1'b0; \
	platform_green_alpha[19][93] = 1'b0; \
	platform_green_alpha[19][94] = 1'b0; \
	platform_green_alpha[19][95] = 1'b1; \
	platform_green_alpha[19][96] = 1'b1; \
	platform_green_alpha[19][97] = 1'b1; \
	platform_green_alpha[19][98] = 1'b1; \
	platform_green_alpha[19][99] = 1'b1; \
	platform_green_alpha[20][0] = 1'b1; \
	platform_green_alpha[20][1] = 1'b1; \
	platform_green_alpha[20][2] = 1'b1; \
	platform_green_alpha[20][3] = 1'b1; \
	platform_green_alpha[20][4] = 1'b1; \
	platform_green_alpha[20][5] = 1'b1; \
	platform_green_alpha[20][6] = 1'b1; \
	platform_green_alpha[20][7] = 1'b1; \
	platform_green_alpha[20][8] = 1'b1; \
	platform_green_alpha[20][9] = 1'b0; \
	platform_green_alpha[20][10] = 1'b0; \
	platform_green_alpha[20][11] = 1'b0; \
	platform_green_alpha[20][12] = 1'b0; \
	platform_green_alpha[20][13] = 1'b0; \
	platform_green_alpha[20][14] = 1'b0; \
	platform_green_alpha[20][15] = 1'b0; \
	platform_green_alpha[20][16] = 1'b0; \
	platform_green_alpha[20][17] = 1'b0; \
	platform_green_alpha[20][18] = 1'b0; \
	platform_green_alpha[20][19] = 1'b0; \
	platform_green_alpha[20][20] = 1'b0; \
	platform_green_alpha[20][21] = 1'b0; \
	platform_green_alpha[20][22] = 1'b0; \
	platform_green_alpha[20][23] = 1'b0; \
	platform_green_alpha[20][24] = 1'b0; \
	platform_green_alpha[20][25] = 1'b0; \
	platform_green_alpha[20][26] = 1'b0; \
	platform_green_alpha[20][27] = 1'b0; \
	platform_green_alpha[20][28] = 1'b0; \
	platform_green_alpha[20][29] = 1'b0; \
	platform_green_alpha[20][30] = 1'b0; \
	platform_green_alpha[20][31] = 1'b0; \
	platform_green_alpha[20][32] = 1'b0; \
	platform_green_alpha[20][33] = 1'b0; \
	platform_green_alpha[20][34] = 1'b0; \
	platform_green_alpha[20][35] = 1'b0; \
	platform_green_alpha[20][36] = 1'b0; \
	platform_green_alpha[20][37] = 1'b0; \
	platform_green_alpha[20][38] = 1'b0; \
	platform_green_alpha[20][39] = 1'b0; \
	platform_green_alpha[20][40] = 1'b0; \
	platform_green_alpha[20][41] = 1'b0; \
	platform_green_alpha[20][42] = 1'b0; \
	platform_green_alpha[20][43] = 1'b0; \
	platform_green_alpha[20][44] = 1'b0; \
	platform_green_alpha[20][45] = 1'b0; \
	platform_green_alpha[20][46] = 1'b0; \
	platform_green_alpha[20][47] = 1'b0; \
	platform_green_alpha[20][48] = 1'b0; \
	platform_green_alpha[20][49] = 1'b0; \
	platform_green_alpha[20][50] = 1'b0; \
	platform_green_alpha[20][51] = 1'b0; \
	platform_green_alpha[20][52] = 1'b0; \
	platform_green_alpha[20][53] = 1'b0; \
	platform_green_alpha[20][54] = 1'b0; \
	platform_green_alpha[20][55] = 1'b0; \
	platform_green_alpha[20][56] = 1'b0; \
	platform_green_alpha[20][57] = 1'b0; \
	platform_green_alpha[20][58] = 1'b0; \
	platform_green_alpha[20][59] = 1'b0; \
	platform_green_alpha[20][60] = 1'b0; \
	platform_green_alpha[20][61] = 1'b0; \
	platform_green_alpha[20][62] = 1'b0; \
	platform_green_alpha[20][63] = 1'b0; \
	platform_green_alpha[20][64] = 1'b0; \
	platform_green_alpha[20][65] = 1'b0; \
	platform_green_alpha[20][66] = 1'b0; \
	platform_green_alpha[20][67] = 1'b0; \
	platform_green_alpha[20][68] = 1'b0; \
	platform_green_alpha[20][69] = 1'b0; \
	platform_green_alpha[20][70] = 1'b0; \
	platform_green_alpha[20][71] = 1'b0; \
	platform_green_alpha[20][72] = 1'b0; \
	platform_green_alpha[20][73] = 1'b0; \
	platform_green_alpha[20][74] = 1'b0; \
	platform_green_alpha[20][75] = 1'b0; \
	platform_green_alpha[20][76] = 1'b0; \
	platform_green_alpha[20][77] = 1'b0; \
	platform_green_alpha[20][78] = 1'b0; \
	platform_green_alpha[20][79] = 1'b0; \
	platform_green_alpha[20][80] = 1'b0; \
	platform_green_alpha[20][81] = 1'b0; \
	platform_green_alpha[20][82] = 1'b0; \
	platform_green_alpha[20][83] = 1'b0; \
	platform_green_alpha[20][84] = 1'b0; \
	platform_green_alpha[20][85] = 1'b0; \
	platform_green_alpha[20][86] = 1'b0; \
	platform_green_alpha[20][87] = 1'b0; \
	platform_green_alpha[20][88] = 1'b0; \
	platform_green_alpha[20][89] = 1'b0; \
	platform_green_alpha[20][90] = 1'b1; \
	platform_green_alpha[20][91] = 1'b1; \
	platform_green_alpha[20][92] = 1'b1; \
	platform_green_alpha[20][93] = 1'b1; \
	platform_green_alpha[20][94] = 1'b1; \
	platform_green_alpha[20][95] = 1'b1; \
	platform_green_alpha[20][96] = 1'b1; \
	platform_green_alpha[20][97] = 1'b1; \
	platform_green_alpha[20][98] = 1'b1; \
	platform_green_alpha[20][99] = 1'b1; \
	platform_green_alpha[21][0] = 1'b1; \
	platform_green_alpha[21][1] = 1'b1; \
	platform_green_alpha[21][2] = 1'b1; \
	platform_green_alpha[21][3] = 1'b1; \
	platform_green_alpha[21][4] = 1'b1; \
	platform_green_alpha[21][5] = 1'b1; \
	platform_green_alpha[21][6] = 1'b1; \
	platform_green_alpha[21][7] = 1'b1; \
	platform_green_alpha[21][8] = 1'b1; \
	platform_green_alpha[21][9] = 1'b0; \
	platform_green_alpha[21][10] = 1'b0; \
	platform_green_alpha[21][11] = 1'b0; \
	platform_green_alpha[21][12] = 1'b0; \
	platform_green_alpha[21][13] = 1'b0; \
	platform_green_alpha[21][14] = 1'b0; \
	platform_green_alpha[21][15] = 1'b0; \
	platform_green_alpha[21][16] = 1'b0; \
	platform_green_alpha[21][17] = 1'b0; \
	platform_green_alpha[21][18] = 1'b0; \
	platform_green_alpha[21][19] = 1'b0; \
	platform_green_alpha[21][20] = 1'b0; \
	platform_green_alpha[21][21] = 1'b0; \
	platform_green_alpha[21][22] = 1'b0; \
	platform_green_alpha[21][23] = 1'b0; \
	platform_green_alpha[21][24] = 1'b0; \
	platform_green_alpha[21][25] = 1'b0; \
	platform_green_alpha[21][26] = 1'b0; \
	platform_green_alpha[21][27] = 1'b0; \
	platform_green_alpha[21][28] = 1'b0; \
	platform_green_alpha[21][29] = 1'b0; \
	platform_green_alpha[21][30] = 1'b0; \
	platform_green_alpha[21][31] = 1'b0; \
	platform_green_alpha[21][32] = 1'b0; \
	platform_green_alpha[21][33] = 1'b0; \
	platform_green_alpha[21][34] = 1'b0; \
	platform_green_alpha[21][35] = 1'b0; \
	platform_green_alpha[21][36] = 1'b0; \
	platform_green_alpha[21][37] = 1'b0; \
	platform_green_alpha[21][38] = 1'b0; \
	platform_green_alpha[21][39] = 1'b0; \
	platform_green_alpha[21][40] = 1'b0; \
	platform_green_alpha[21][41] = 1'b0; \
	platform_green_alpha[21][42] = 1'b0; \
	platform_green_alpha[21][43] = 1'b0; \
	platform_green_alpha[21][44] = 1'b0; \
	platform_green_alpha[21][45] = 1'b0; \
	platform_green_alpha[21][46] = 1'b0; \
	platform_green_alpha[21][47] = 1'b0; \
	platform_green_alpha[21][48] = 1'b0; \
	platform_green_alpha[21][49] = 1'b0; \
	platform_green_alpha[21][50] = 1'b0; \
	platform_green_alpha[21][51] = 1'b0; \
	platform_green_alpha[21][52] = 1'b0; \
	platform_green_alpha[21][53] = 1'b0; \
	platform_green_alpha[21][54] = 1'b0; \
	platform_green_alpha[21][55] = 1'b0; \
	platform_green_alpha[21][56] = 1'b0; \
	platform_green_alpha[21][57] = 1'b0; \
	platform_green_alpha[21][58] = 1'b0; \
	platform_green_alpha[21][59] = 1'b0; \
	platform_green_alpha[21][60] = 1'b0; \
	platform_green_alpha[21][61] = 1'b0; \
	platform_green_alpha[21][62] = 1'b0; \
	platform_green_alpha[21][63] = 1'b0; \
	platform_green_alpha[21][64] = 1'b0; \
	platform_green_alpha[21][65] = 1'b0; \
	platform_green_alpha[21][66] = 1'b0; \
	platform_green_alpha[21][67] = 1'b0; \
	platform_green_alpha[21][68] = 1'b0; \
	platform_green_alpha[21][69] = 1'b0; \
	platform_green_alpha[21][70] = 1'b0; \
	platform_green_alpha[21][71] = 1'b0; \
	platform_green_alpha[21][72] = 1'b0; \
	platform_green_alpha[21][73] = 1'b0; \
	platform_green_alpha[21][74] = 1'b0; \
	platform_green_alpha[21][75] = 1'b0; \
	platform_green_alpha[21][76] = 1'b0; \
	platform_green_alpha[21][77] = 1'b0; \
	platform_green_alpha[21][78] = 1'b0; \
	platform_green_alpha[21][79] = 1'b0; \
	platform_green_alpha[21][80] = 1'b0; \
	platform_green_alpha[21][81] = 1'b0; \
	platform_green_alpha[21][82] = 1'b0; \
	platform_green_alpha[21][83] = 1'b0; \
	platform_green_alpha[21][84] = 1'b0; \
	platform_green_alpha[21][85] = 1'b0; \
	platform_green_alpha[21][86] = 1'b0; \
	platform_green_alpha[21][87] = 1'b0; \
	platform_green_alpha[21][88] = 1'b0; \
	platform_green_alpha[21][89] = 1'b0; \
	platform_green_alpha[21][90] = 1'b1; \
	platform_green_alpha[21][91] = 1'b1; \
	platform_green_alpha[21][92] = 1'b1; \
	platform_green_alpha[21][93] = 1'b1; \
	platform_green_alpha[21][94] = 1'b1; \
	platform_green_alpha[21][95] = 1'b1; \
	platform_green_alpha[21][96] = 1'b1; \
	platform_green_alpha[21][97] = 1'b1; \
	platform_green_alpha[21][98] = 1'b1; \
	platform_green_alpha[21][99] = 1'b1; \
	platform_green_alpha[22][0] = 1'b1; \
	platform_green_alpha[22][1] = 1'b1; \
	platform_green_alpha[22][2] = 1'b1; \
	platform_green_alpha[22][3] = 1'b1; \
	platform_green_alpha[22][4] = 1'b1; \
	platform_green_alpha[22][5] = 1'b1; \
	platform_green_alpha[22][6] = 1'b1; \
	platform_green_alpha[22][7] = 1'b1; \
	platform_green_alpha[22][8] = 1'b1; \
	platform_green_alpha[22][9] = 1'b0; \
	platform_green_alpha[22][10] = 1'b0; \
	platform_green_alpha[22][11] = 1'b0; \
	platform_green_alpha[22][12] = 1'b0; \
	platform_green_alpha[22][13] = 1'b0; \
	platform_green_alpha[22][14] = 1'b0; \
	platform_green_alpha[22][15] = 1'b0; \
	platform_green_alpha[22][16] = 1'b0; \
	platform_green_alpha[22][17] = 1'b0; \
	platform_green_alpha[22][18] = 1'b0; \
	platform_green_alpha[22][19] = 1'b0; \
	platform_green_alpha[22][20] = 1'b0; \
	platform_green_alpha[22][21] = 1'b0; \
	platform_green_alpha[22][22] = 1'b0; \
	platform_green_alpha[22][23] = 1'b0; \
	platform_green_alpha[22][24] = 1'b0; \
	platform_green_alpha[22][25] = 1'b0; \
	platform_green_alpha[22][26] = 1'b0; \
	platform_green_alpha[22][27] = 1'b0; \
	platform_green_alpha[22][28] = 1'b0; \
	platform_green_alpha[22][29] = 1'b0; \
	platform_green_alpha[22][30] = 1'b0; \
	platform_green_alpha[22][31] = 1'b0; \
	platform_green_alpha[22][32] = 1'b0; \
	platform_green_alpha[22][33] = 1'b0; \
	platform_green_alpha[22][34] = 1'b0; \
	platform_green_alpha[22][35] = 1'b0; \
	platform_green_alpha[22][36] = 1'b0; \
	platform_green_alpha[22][37] = 1'b0; \
	platform_green_alpha[22][38] = 1'b0; \
	platform_green_alpha[22][39] = 1'b0; \
	platform_green_alpha[22][40] = 1'b0; \
	platform_green_alpha[22][41] = 1'b0; \
	platform_green_alpha[22][42] = 1'b0; \
	platform_green_alpha[22][43] = 1'b0; \
	platform_green_alpha[22][44] = 1'b0; \
	platform_green_alpha[22][45] = 1'b0; \
	platform_green_alpha[22][46] = 1'b0; \
	platform_green_alpha[22][47] = 1'b0; \
	platform_green_alpha[22][48] = 1'b0; \
	platform_green_alpha[22][49] = 1'b0; \
	platform_green_alpha[22][50] = 1'b0; \
	platform_green_alpha[22][51] = 1'b0; \
	platform_green_alpha[22][52] = 1'b0; \
	platform_green_alpha[22][53] = 1'b0; \
	platform_green_alpha[22][54] = 1'b0; \
	platform_green_alpha[22][55] = 1'b0; \
	platform_green_alpha[22][56] = 1'b0; \
	platform_green_alpha[22][57] = 1'b0; \
	platform_green_alpha[22][58] = 1'b0; \
	platform_green_alpha[22][59] = 1'b0; \
	platform_green_alpha[22][60] = 1'b0; \
	platform_green_alpha[22][61] = 1'b0; \
	platform_green_alpha[22][62] = 1'b0; \
	platform_green_alpha[22][63] = 1'b0; \
	platform_green_alpha[22][64] = 1'b0; \
	platform_green_alpha[22][65] = 1'b0; \
	platform_green_alpha[22][66] = 1'b0; \
	platform_green_alpha[22][67] = 1'b0; \
	platform_green_alpha[22][68] = 1'b0; \
	platform_green_alpha[22][69] = 1'b0; \
	platform_green_alpha[22][70] = 1'b0; \
	platform_green_alpha[22][71] = 1'b0; \
	platform_green_alpha[22][72] = 1'b0; \
	platform_green_alpha[22][73] = 1'b0; \
	platform_green_alpha[22][74] = 1'b0; \
	platform_green_alpha[22][75] = 1'b0; \
	platform_green_alpha[22][76] = 1'b0; \
	platform_green_alpha[22][77] = 1'b0; \
	platform_green_alpha[22][78] = 1'b0; \
	platform_green_alpha[22][79] = 1'b0; \
	platform_green_alpha[22][80] = 1'b0; \
	platform_green_alpha[22][81] = 1'b0; \
	platform_green_alpha[22][82] = 1'b0; \
	platform_green_alpha[22][83] = 1'b0; \
	platform_green_alpha[22][84] = 1'b0; \
	platform_green_alpha[22][85] = 1'b0; \
	platform_green_alpha[22][86] = 1'b0; \
	platform_green_alpha[22][87] = 1'b0; \
	platform_green_alpha[22][88] = 1'b0; \
	platform_green_alpha[22][89] = 1'b0; \
	platform_green_alpha[22][90] = 1'b1; \
	platform_green_alpha[22][91] = 1'b1; \
	platform_green_alpha[22][92] = 1'b1; \
	platform_green_alpha[22][93] = 1'b1; \
	platform_green_alpha[22][94] = 1'b1; \
	platform_green_alpha[22][95] = 1'b1; \
	platform_green_alpha[22][96] = 1'b1; \
	platform_green_alpha[22][97] = 1'b1; \
	platform_green_alpha[22][98] = 1'b1; \
	platform_green_alpha[22][99] = 1'b1; \
	platform_green_alpha[23][0] = 1'b1; \
	platform_green_alpha[23][1] = 1'b1; \
	platform_green_alpha[23][2] = 1'b1; \
	platform_green_alpha[23][3] = 1'b1; \
	platform_green_alpha[23][4] = 1'b1; \
	platform_green_alpha[23][5] = 1'b1; \
	platform_green_alpha[23][6] = 1'b1; \
	platform_green_alpha[23][7] = 1'b1; \
	platform_green_alpha[23][8] = 1'b1; \
	platform_green_alpha[23][9] = 1'b0; \
	platform_green_alpha[23][10] = 1'b0; \
	platform_green_alpha[23][11] = 1'b0; \
	platform_green_alpha[23][12] = 1'b0; \
	platform_green_alpha[23][13] = 1'b0; \
	platform_green_alpha[23][14] = 1'b0; \
	platform_green_alpha[23][15] = 1'b0; \
	platform_green_alpha[23][16] = 1'b0; \
	platform_green_alpha[23][17] = 1'b0; \
	platform_green_alpha[23][18] = 1'b0; \
	platform_green_alpha[23][19] = 1'b0; \
	platform_green_alpha[23][20] = 1'b0; \
	platform_green_alpha[23][21] = 1'b0; \
	platform_green_alpha[23][22] = 1'b0; \
	platform_green_alpha[23][23] = 1'b0; \
	platform_green_alpha[23][24] = 1'b0; \
	platform_green_alpha[23][25] = 1'b0; \
	platform_green_alpha[23][26] = 1'b0; \
	platform_green_alpha[23][27] = 1'b0; \
	platform_green_alpha[23][28] = 1'b0; \
	platform_green_alpha[23][29] = 1'b0; \
	platform_green_alpha[23][30] = 1'b0; \
	platform_green_alpha[23][31] = 1'b0; \
	platform_green_alpha[23][32] = 1'b0; \
	platform_green_alpha[23][33] = 1'b0; \
	platform_green_alpha[23][34] = 1'b0; \
	platform_green_alpha[23][35] = 1'b0; \
	platform_green_alpha[23][36] = 1'b0; \
	platform_green_alpha[23][37] = 1'b0; \
	platform_green_alpha[23][38] = 1'b0; \
	platform_green_alpha[23][39] = 1'b0; \
	platform_green_alpha[23][40] = 1'b0; \
	platform_green_alpha[23][41] = 1'b0; \
	platform_green_alpha[23][42] = 1'b0; \
	platform_green_alpha[23][43] = 1'b0; \
	platform_green_alpha[23][44] = 1'b0; \
	platform_green_alpha[23][45] = 1'b0; \
	platform_green_alpha[23][46] = 1'b0; \
	platform_green_alpha[23][47] = 1'b0; \
	platform_green_alpha[23][48] = 1'b0; \
	platform_green_alpha[23][49] = 1'b0; \
	platform_green_alpha[23][50] = 1'b0; \
	platform_green_alpha[23][51] = 1'b0; \
	platform_green_alpha[23][52] = 1'b0; \
	platform_green_alpha[23][53] = 1'b0; \
	platform_green_alpha[23][54] = 1'b0; \
	platform_green_alpha[23][55] = 1'b0; \
	platform_green_alpha[23][56] = 1'b0; \
	platform_green_alpha[23][57] = 1'b0; \
	platform_green_alpha[23][58] = 1'b0; \
	platform_green_alpha[23][59] = 1'b0; \
	platform_green_alpha[23][60] = 1'b0; \
	platform_green_alpha[23][61] = 1'b0; \
	platform_green_alpha[23][62] = 1'b0; \
	platform_green_alpha[23][63] = 1'b0; \
	platform_green_alpha[23][64] = 1'b0; \
	platform_green_alpha[23][65] = 1'b0; \
	platform_green_alpha[23][66] = 1'b0; \
	platform_green_alpha[23][67] = 1'b0; \
	platform_green_alpha[23][68] = 1'b0; \
	platform_green_alpha[23][69] = 1'b0; \
	platform_green_alpha[23][70] = 1'b0; \
	platform_green_alpha[23][71] = 1'b0; \
	platform_green_alpha[23][72] = 1'b0; \
	platform_green_alpha[23][73] = 1'b0; \
	platform_green_alpha[23][74] = 1'b0; \
	platform_green_alpha[23][75] = 1'b0; \
	platform_green_alpha[23][76] = 1'b0; \
	platform_green_alpha[23][77] = 1'b0; \
	platform_green_alpha[23][78] = 1'b0; \
	platform_green_alpha[23][79] = 1'b0; \
	platform_green_alpha[23][80] = 1'b0; \
	platform_green_alpha[23][81] = 1'b0; \
	platform_green_alpha[23][82] = 1'b0; \
	platform_green_alpha[23][83] = 1'b0; \
	platform_green_alpha[23][84] = 1'b0; \
	platform_green_alpha[23][85] = 1'b0; \
	platform_green_alpha[23][86] = 1'b0; \
	platform_green_alpha[23][87] = 1'b0; \
	platform_green_alpha[23][88] = 1'b0; \
	platform_green_alpha[23][89] = 1'b0; \
	platform_green_alpha[23][90] = 1'b1; \
	platform_green_alpha[23][91] = 1'b1; \
	platform_green_alpha[23][92] = 1'b1; \
	platform_green_alpha[23][93] = 1'b1; \
	platform_green_alpha[23][94] = 1'b1; \
	platform_green_alpha[23][95] = 1'b1; \
	platform_green_alpha[23][96] = 1'b1; \
	platform_green_alpha[23][97] = 1'b1; \
	platform_green_alpha[23][98] = 1'b1; \
	platform_green_alpha[23][99] = 1'b1; \
	platform_green_alpha[24][0] = 1'b1; \
	platform_green_alpha[24][1] = 1'b1; \
	platform_green_alpha[24][2] = 1'b1; \
	platform_green_alpha[24][3] = 1'b1; \
	platform_green_alpha[24][4] = 1'b1; \
	platform_green_alpha[24][5] = 1'b1; \
	platform_green_alpha[24][6] = 1'b1; \
	platform_green_alpha[24][7] = 1'b1; \
	platform_green_alpha[24][8] = 1'b1; \
	platform_green_alpha[24][9] = 1'b0; \
	platform_green_alpha[24][10] = 1'b0; \
	platform_green_alpha[24][11] = 1'b0; \
	platform_green_alpha[24][12] = 1'b0; \
	platform_green_alpha[24][13] = 1'b0; \
	platform_green_alpha[24][14] = 1'b0; \
	platform_green_alpha[24][15] = 1'b0; \
	platform_green_alpha[24][16] = 1'b0; \
	platform_green_alpha[24][17] = 1'b0; \
	platform_green_alpha[24][18] = 1'b0; \
	platform_green_alpha[24][19] = 1'b0; \
	platform_green_alpha[24][20] = 1'b0; \
	platform_green_alpha[24][21] = 1'b0; \
	platform_green_alpha[24][22] = 1'b0; \
	platform_green_alpha[24][23] = 1'b0; \
	platform_green_alpha[24][24] = 1'b0; \
	platform_green_alpha[24][25] = 1'b0; \
	platform_green_alpha[24][26] = 1'b0; \
	platform_green_alpha[24][27] = 1'b0; \
	platform_green_alpha[24][28] = 1'b0; \
	platform_green_alpha[24][29] = 1'b0; \
	platform_green_alpha[24][30] = 1'b0; \
	platform_green_alpha[24][31] = 1'b0; \
	platform_green_alpha[24][32] = 1'b0; \
	platform_green_alpha[24][33] = 1'b0; \
	platform_green_alpha[24][34] = 1'b0; \
	platform_green_alpha[24][35] = 1'b0; \
	platform_green_alpha[24][36] = 1'b0; \
	platform_green_alpha[24][37] = 1'b0; \
	platform_green_alpha[24][38] = 1'b0; \
	platform_green_alpha[24][39] = 1'b0; \
	platform_green_alpha[24][40] = 1'b0; \
	platform_green_alpha[24][41] = 1'b0; \
	platform_green_alpha[24][42] = 1'b0; \
	platform_green_alpha[24][43] = 1'b0; \
	platform_green_alpha[24][44] = 1'b0; \
	platform_green_alpha[24][45] = 1'b0; \
	platform_green_alpha[24][46] = 1'b0; \
	platform_green_alpha[24][47] = 1'b0; \
	platform_green_alpha[24][48] = 1'b0; \
	platform_green_alpha[24][49] = 1'b0; \
	platform_green_alpha[24][50] = 1'b0; \
	platform_green_alpha[24][51] = 1'b0; \
	platform_green_alpha[24][52] = 1'b0; \
	platform_green_alpha[24][53] = 1'b0; \
	platform_green_alpha[24][54] = 1'b0; \
	platform_green_alpha[24][55] = 1'b0; \
	platform_green_alpha[24][56] = 1'b0; \
	platform_green_alpha[24][57] = 1'b0; \
	platform_green_alpha[24][58] = 1'b0; \
	platform_green_alpha[24][59] = 1'b0; \
	platform_green_alpha[24][60] = 1'b0; \
	platform_green_alpha[24][61] = 1'b0; \
	platform_green_alpha[24][62] = 1'b0; \
	platform_green_alpha[24][63] = 1'b0; \
	platform_green_alpha[24][64] = 1'b0; \
	platform_green_alpha[24][65] = 1'b0; \
	platform_green_alpha[24][66] = 1'b0; \
	platform_green_alpha[24][67] = 1'b0; \
	platform_green_alpha[24][68] = 1'b0; \
	platform_green_alpha[24][69] = 1'b0; \
	platform_green_alpha[24][70] = 1'b0; \
	platform_green_alpha[24][71] = 1'b0; \
	platform_green_alpha[24][72] = 1'b0; \
	platform_green_alpha[24][73] = 1'b0; \
	platform_green_alpha[24][74] = 1'b0; \
	platform_green_alpha[24][75] = 1'b0; \
	platform_green_alpha[24][76] = 1'b0; \
	platform_green_alpha[24][77] = 1'b0; \
	platform_green_alpha[24][78] = 1'b0; \
	platform_green_alpha[24][79] = 1'b0; \
	platform_green_alpha[24][80] = 1'b0; \
	platform_green_alpha[24][81] = 1'b0; \
	platform_green_alpha[24][82] = 1'b0; \
	platform_green_alpha[24][83] = 1'b0; \
	platform_green_alpha[24][84] = 1'b0; \
	platform_green_alpha[24][85] = 1'b0; \
	platform_green_alpha[24][86] = 1'b0; \
	platform_green_alpha[24][87] = 1'b0; \
	platform_green_alpha[24][88] = 1'b0; \
	platform_green_alpha[24][89] = 1'b0; \
	platform_green_alpha[24][90] = 1'b1; \
	platform_green_alpha[24][91] = 1'b1; \
	platform_green_alpha[24][92] = 1'b1; \
	platform_green_alpha[24][93] = 1'b1; \
	platform_green_alpha[24][94] = 1'b1; \
	platform_green_alpha[24][95] = 1'b1; \
	platform_green_alpha[24][96] = 1'b1; \
	platform_green_alpha[24][97] = 1'b1; \
	platform_green_alpha[24][98] = 1'b1; \
	platform_green_alpha[24][99] = 1'b1; \
	platform_green_alpha[25][0] = 1'b1; \
	platform_green_alpha[25][1] = 1'b1; \
	platform_green_alpha[25][2] = 1'b1; \
	platform_green_alpha[25][3] = 1'b1; \
	platform_green_alpha[25][4] = 1'b1; \
	platform_green_alpha[25][5] = 1'b1; \
	platform_green_alpha[25][6] = 1'b1; \
	platform_green_alpha[25][7] = 1'b1; \
	platform_green_alpha[25][8] = 1'b1; \
	platform_green_alpha[25][9] = 1'b1; \
	platform_green_alpha[25][10] = 1'b1; \
	platform_green_alpha[25][11] = 1'b1; \
	platform_green_alpha[25][12] = 1'b1; \
	platform_green_alpha[25][13] = 1'b1; \
	platform_green_alpha[25][14] = 1'b1; \
	platform_green_alpha[25][15] = 1'b1; \
	platform_green_alpha[25][16] = 1'b1; \
	platform_green_alpha[25][17] = 1'b1; \
	platform_green_alpha[25][18] = 1'b1; \
	platform_green_alpha[25][19] = 1'b1; \
	platform_green_alpha[25][20] = 1'b1; \
	platform_green_alpha[25][21] = 1'b1; \
	platform_green_alpha[25][22] = 1'b1; \
	platform_green_alpha[25][23] = 1'b1; \
	platform_green_alpha[25][24] = 1'b1; \
	platform_green_alpha[25][25] = 1'b1; \
	platform_green_alpha[25][26] = 1'b1; \
	platform_green_alpha[25][27] = 1'b1; \
	platform_green_alpha[25][28] = 1'b1; \
	platform_green_alpha[25][29] = 1'b1; \
	platform_green_alpha[25][30] = 1'b1; \
	platform_green_alpha[25][31] = 1'b1; \
	platform_green_alpha[25][32] = 1'b1; \
	platform_green_alpha[25][33] = 1'b1; \
	platform_green_alpha[25][34] = 1'b1; \
	platform_green_alpha[25][35] = 1'b1; \
	platform_green_alpha[25][36] = 1'b1; \
	platform_green_alpha[25][37] = 1'b1; \
	platform_green_alpha[25][38] = 1'b1; \
	platform_green_alpha[25][39] = 1'b1; \
	platform_green_alpha[25][40] = 1'b1; \
	platform_green_alpha[25][41] = 1'b1; \
	platform_green_alpha[25][42] = 1'b1; \
	platform_green_alpha[25][43] = 1'b1; \
	platform_green_alpha[25][44] = 1'b1; \
	platform_green_alpha[25][45] = 1'b1; \
	platform_green_alpha[25][46] = 1'b1; \
	platform_green_alpha[25][47] = 1'b1; \
	platform_green_alpha[25][48] = 1'b1; \
	platform_green_alpha[25][49] = 1'b1; \
	platform_green_alpha[25][50] = 1'b1; \
	platform_green_alpha[25][51] = 1'b1; \
	platform_green_alpha[25][52] = 1'b1; \
	platform_green_alpha[25][53] = 1'b1; \
	platform_green_alpha[25][54] = 1'b1; \
	platform_green_alpha[25][55] = 1'b1; \
	platform_green_alpha[25][56] = 1'b1; \
	platform_green_alpha[25][57] = 1'b1; \
	platform_green_alpha[25][58] = 1'b1; \
	platform_green_alpha[25][59] = 1'b1; \
	platform_green_alpha[25][60] = 1'b1; \
	platform_green_alpha[25][61] = 1'b1; \
	platform_green_alpha[25][62] = 1'b1; \
	platform_green_alpha[25][63] = 1'b1; \
	platform_green_alpha[25][64] = 1'b1; \
	platform_green_alpha[25][65] = 1'b1; \
	platform_green_alpha[25][66] = 1'b1; \
	platform_green_alpha[25][67] = 1'b1; \
	platform_green_alpha[25][68] = 1'b1; \
	platform_green_alpha[25][69] = 1'b1; \
	platform_green_alpha[25][70] = 1'b1; \
	platform_green_alpha[25][71] = 1'b1; \
	platform_green_alpha[25][72] = 1'b1; \
	platform_green_alpha[25][73] = 1'b1; \
	platform_green_alpha[25][74] = 1'b1; \
	platform_green_alpha[25][75] = 1'b1; \
	platform_green_alpha[25][76] = 1'b1; \
	platform_green_alpha[25][77] = 1'b1; \
	platform_green_alpha[25][78] = 1'b1; \
	platform_green_alpha[25][79] = 1'b1; \
	platform_green_alpha[25][80] = 1'b1; \
	platform_green_alpha[25][81] = 1'b1; \
	platform_green_alpha[25][82] = 1'b1; \
	platform_green_alpha[25][83] = 1'b1; \
	platform_green_alpha[25][84] = 1'b1; \
	platform_green_alpha[25][85] = 1'b1; \
	platform_green_alpha[25][86] = 1'b1; \
	platform_green_alpha[25][87] = 1'b1; \
	platform_green_alpha[25][88] = 1'b1; \
	platform_green_alpha[25][89] = 1'b1; \
	platform_green_alpha[25][90] = 1'b1; \
	platform_green_alpha[25][91] = 1'b1; \
	platform_green_alpha[25][92] = 1'b1; \
	platform_green_alpha[25][93] = 1'b1; \
	platform_green_alpha[25][94] = 1'b1; \
	platform_green_alpha[25][95] = 1'b1; \
	platform_green_alpha[25][96] = 1'b1; \
	platform_green_alpha[25][97] = 1'b1; \
	platform_green_alpha[25][98] = 1'b1; \
	platform_green_alpha[25][99] = 1'b1; \
	platform_green_alpha[26][0] = 1'b1; \
	platform_green_alpha[26][1] = 1'b1; \
	platform_green_alpha[26][2] = 1'b1; \
	platform_green_alpha[26][3] = 1'b1; \
	platform_green_alpha[26][4] = 1'b1; \
	platform_green_alpha[26][5] = 1'b1; \
	platform_green_alpha[26][6] = 1'b1; \
	platform_green_alpha[26][7] = 1'b1; \
	platform_green_alpha[26][8] = 1'b1; \
	platform_green_alpha[26][9] = 1'b1; \
	platform_green_alpha[26][10] = 1'b1; \
	platform_green_alpha[26][11] = 1'b1; \
	platform_green_alpha[26][12] = 1'b1; \
	platform_green_alpha[26][13] = 1'b1; \
	platform_green_alpha[26][14] = 1'b1; \
	platform_green_alpha[26][15] = 1'b1; \
	platform_green_alpha[26][16] = 1'b1; \
	platform_green_alpha[26][17] = 1'b1; \
	platform_green_alpha[26][18] = 1'b1; \
	platform_green_alpha[26][19] = 1'b1; \
	platform_green_alpha[26][20] = 1'b1; \
	platform_green_alpha[26][21] = 1'b1; \
	platform_green_alpha[26][22] = 1'b1; \
	platform_green_alpha[26][23] = 1'b1; \
	platform_green_alpha[26][24] = 1'b1; \
	platform_green_alpha[26][25] = 1'b1; \
	platform_green_alpha[26][26] = 1'b1; \
	platform_green_alpha[26][27] = 1'b1; \
	platform_green_alpha[26][28] = 1'b1; \
	platform_green_alpha[26][29] = 1'b1; \
	platform_green_alpha[26][30] = 1'b1; \
	platform_green_alpha[26][31] = 1'b1; \
	platform_green_alpha[26][32] = 1'b1; \
	platform_green_alpha[26][33] = 1'b1; \
	platform_green_alpha[26][34] = 1'b1; \
	platform_green_alpha[26][35] = 1'b1; \
	platform_green_alpha[26][36] = 1'b1; \
	platform_green_alpha[26][37] = 1'b1; \
	platform_green_alpha[26][38] = 1'b1; \
	platform_green_alpha[26][39] = 1'b1; \
	platform_green_alpha[26][40] = 1'b1; \
	platform_green_alpha[26][41] = 1'b1; \
	platform_green_alpha[26][42] = 1'b1; \
	platform_green_alpha[26][43] = 1'b1; \
	platform_green_alpha[26][44] = 1'b1; \
	platform_green_alpha[26][45] = 1'b1; \
	platform_green_alpha[26][46] = 1'b1; \
	platform_green_alpha[26][47] = 1'b1; \
	platform_green_alpha[26][48] = 1'b1; \
	platform_green_alpha[26][49] = 1'b1; \
	platform_green_alpha[26][50] = 1'b1; \
	platform_green_alpha[26][51] = 1'b1; \
	platform_green_alpha[26][52] = 1'b1; \
	platform_green_alpha[26][53] = 1'b1; \
	platform_green_alpha[26][54] = 1'b1; \
	platform_green_alpha[26][55] = 1'b1; \
	platform_green_alpha[26][56] = 1'b1; \
	platform_green_alpha[26][57] = 1'b1; \
	platform_green_alpha[26][58] = 1'b1; \
	platform_green_alpha[26][59] = 1'b1; \
	platform_green_alpha[26][60] = 1'b1; \
	platform_green_alpha[26][61] = 1'b1; \
	platform_green_alpha[26][62] = 1'b1; \
	platform_green_alpha[26][63] = 1'b1; \
	platform_green_alpha[26][64] = 1'b1; \
	platform_green_alpha[26][65] = 1'b1; \
	platform_green_alpha[26][66] = 1'b1; \
	platform_green_alpha[26][67] = 1'b1; \
	platform_green_alpha[26][68] = 1'b1; \
	platform_green_alpha[26][69] = 1'b1; \
	platform_green_alpha[26][70] = 1'b1; \
	platform_green_alpha[26][71] = 1'b1; \
	platform_green_alpha[26][72] = 1'b1; \
	platform_green_alpha[26][73] = 1'b1; \
	platform_green_alpha[26][74] = 1'b1; \
	platform_green_alpha[26][75] = 1'b1; \
	platform_green_alpha[26][76] = 1'b1; \
	platform_green_alpha[26][77] = 1'b1; \
	platform_green_alpha[26][78] = 1'b1; \
	platform_green_alpha[26][79] = 1'b1; \
	platform_green_alpha[26][80] = 1'b1; \
	platform_green_alpha[26][81] = 1'b1; \
	platform_green_alpha[26][82] = 1'b1; \
	platform_green_alpha[26][83] = 1'b1; \
	platform_green_alpha[26][84] = 1'b1; \
	platform_green_alpha[26][85] = 1'b1; \
	platform_green_alpha[26][86] = 1'b1; \
	platform_green_alpha[26][87] = 1'b1; \
	platform_green_alpha[26][88] = 1'b1; \
	platform_green_alpha[26][89] = 1'b1; \
	platform_green_alpha[26][90] = 1'b1; \
	platform_green_alpha[26][91] = 1'b1; \
	platform_green_alpha[26][92] = 1'b1; \
	platform_green_alpha[26][93] = 1'b1; \
	platform_green_alpha[26][94] = 1'b1; \
	platform_green_alpha[26][95] = 1'b1; \
	platform_green_alpha[26][96] = 1'b1; \
	platform_green_alpha[26][97] = 1'b1; \
	platform_green_alpha[26][98] = 1'b1; \
	platform_green_alpha[26][99] = 1'b1; \
	platform_green_alpha[27][0] = 1'b1; \
	platform_green_alpha[27][1] = 1'b1; \
	platform_green_alpha[27][2] = 1'b1; \
	platform_green_alpha[27][3] = 1'b1; \
	platform_green_alpha[27][4] = 1'b1; \
	platform_green_alpha[27][5] = 1'b1; \
	platform_green_alpha[27][6] = 1'b1; \
	platform_green_alpha[27][7] = 1'b1; \
	platform_green_alpha[27][8] = 1'b1; \
	platform_green_alpha[27][9] = 1'b1; \
	platform_green_alpha[27][10] = 1'b1; \
	platform_green_alpha[27][11] = 1'b1; \
	platform_green_alpha[27][12] = 1'b1; \
	platform_green_alpha[27][13] = 1'b1; \
	platform_green_alpha[27][14] = 1'b1; \
	platform_green_alpha[27][15] = 1'b1; \
	platform_green_alpha[27][16] = 1'b1; \
	platform_green_alpha[27][17] = 1'b1; \
	platform_green_alpha[27][18] = 1'b1; \
	platform_green_alpha[27][19] = 1'b1; \
	platform_green_alpha[27][20] = 1'b1; \
	platform_green_alpha[27][21] = 1'b1; \
	platform_green_alpha[27][22] = 1'b1; \
	platform_green_alpha[27][23] = 1'b1; \
	platform_green_alpha[27][24] = 1'b1; \
	platform_green_alpha[27][25] = 1'b1; \
	platform_green_alpha[27][26] = 1'b1; \
	platform_green_alpha[27][27] = 1'b1; \
	platform_green_alpha[27][28] = 1'b1; \
	platform_green_alpha[27][29] = 1'b1; \
	platform_green_alpha[27][30] = 1'b1; \
	platform_green_alpha[27][31] = 1'b1; \
	platform_green_alpha[27][32] = 1'b1; \
	platform_green_alpha[27][33] = 1'b1; \
	platform_green_alpha[27][34] = 1'b1; \
	platform_green_alpha[27][35] = 1'b1; \
	platform_green_alpha[27][36] = 1'b1; \
	platform_green_alpha[27][37] = 1'b1; \
	platform_green_alpha[27][38] = 1'b1; \
	platform_green_alpha[27][39] = 1'b1; \
	platform_green_alpha[27][40] = 1'b1; \
	platform_green_alpha[27][41] = 1'b1; \
	platform_green_alpha[27][42] = 1'b1; \
	platform_green_alpha[27][43] = 1'b1; \
	platform_green_alpha[27][44] = 1'b1; \
	platform_green_alpha[27][45] = 1'b1; \
	platform_green_alpha[27][46] = 1'b1; \
	platform_green_alpha[27][47] = 1'b1; \
	platform_green_alpha[27][48] = 1'b1; \
	platform_green_alpha[27][49] = 1'b1; \
	platform_green_alpha[27][50] = 1'b1; \
	platform_green_alpha[27][51] = 1'b1; \
	platform_green_alpha[27][52] = 1'b1; \
	platform_green_alpha[27][53] = 1'b1; \
	platform_green_alpha[27][54] = 1'b1; \
	platform_green_alpha[27][55] = 1'b1; \
	platform_green_alpha[27][56] = 1'b1; \
	platform_green_alpha[27][57] = 1'b1; \
	platform_green_alpha[27][58] = 1'b1; \
	platform_green_alpha[27][59] = 1'b1; \
	platform_green_alpha[27][60] = 1'b1; \
	platform_green_alpha[27][61] = 1'b1; \
	platform_green_alpha[27][62] = 1'b1; \
	platform_green_alpha[27][63] = 1'b1; \
	platform_green_alpha[27][64] = 1'b1; \
	platform_green_alpha[27][65] = 1'b1; \
	platform_green_alpha[27][66] = 1'b1; \
	platform_green_alpha[27][67] = 1'b1; \
	platform_green_alpha[27][68] = 1'b1; \
	platform_green_alpha[27][69] = 1'b1; \
	platform_green_alpha[27][70] = 1'b1; \
	platform_green_alpha[27][71] = 1'b1; \
	platform_green_alpha[27][72] = 1'b1; \
	platform_green_alpha[27][73] = 1'b1; \
	platform_green_alpha[27][74] = 1'b1; \
	platform_green_alpha[27][75] = 1'b1; \
	platform_green_alpha[27][76] = 1'b1; \
	platform_green_alpha[27][77] = 1'b1; \
	platform_green_alpha[27][78] = 1'b1; \
	platform_green_alpha[27][79] = 1'b1; \
	platform_green_alpha[27][80] = 1'b1; \
	platform_green_alpha[27][81] = 1'b1; \
	platform_green_alpha[27][82] = 1'b1; \
	platform_green_alpha[27][83] = 1'b1; \
	platform_green_alpha[27][84] = 1'b1; \
	platform_green_alpha[27][85] = 1'b1; \
	platform_green_alpha[27][86] = 1'b1; \
	platform_green_alpha[27][87] = 1'b1; \
	platform_green_alpha[27][88] = 1'b1; \
	platform_green_alpha[27][89] = 1'b1; \
	platform_green_alpha[27][90] = 1'b1; \
	platform_green_alpha[27][91] = 1'b1; \
	platform_green_alpha[27][92] = 1'b1; \
	platform_green_alpha[27][93] = 1'b1; \
	platform_green_alpha[27][94] = 1'b1; \
	platform_green_alpha[27][95] = 1'b1; \
	platform_green_alpha[27][96] = 1'b1; \
	platform_green_alpha[27][97] = 1'b1; \
	platform_green_alpha[27][98] = 1'b1; \
	platform_green_alpha[27][99] = 1'b1; \
	platform_green_alpha[28][0] = 1'b1; \
	platform_green_alpha[28][1] = 1'b1; \
	platform_green_alpha[28][2] = 1'b1; \
	platform_green_alpha[28][3] = 1'b1; \
	platform_green_alpha[28][4] = 1'b1; \
	platform_green_alpha[28][5] = 1'b1; \
	platform_green_alpha[28][6] = 1'b1; \
	platform_green_alpha[28][7] = 1'b1; \
	platform_green_alpha[28][8] = 1'b1; \
	platform_green_alpha[28][9] = 1'b1; \
	platform_green_alpha[28][10] = 1'b1; \
	platform_green_alpha[28][11] = 1'b1; \
	platform_green_alpha[28][12] = 1'b1; \
	platform_green_alpha[28][13] = 1'b1; \
	platform_green_alpha[28][14] = 1'b1; \
	platform_green_alpha[28][15] = 1'b1; \
	platform_green_alpha[28][16] = 1'b1; \
	platform_green_alpha[28][17] = 1'b1; \
	platform_green_alpha[28][18] = 1'b1; \
	platform_green_alpha[28][19] = 1'b1; \
	platform_green_alpha[28][20] = 1'b1; \
	platform_green_alpha[28][21] = 1'b1; \
	platform_green_alpha[28][22] = 1'b1; \
	platform_green_alpha[28][23] = 1'b1; \
	platform_green_alpha[28][24] = 1'b1; \
	platform_green_alpha[28][25] = 1'b1; \
	platform_green_alpha[28][26] = 1'b1; \
	platform_green_alpha[28][27] = 1'b1; \
	platform_green_alpha[28][28] = 1'b1; \
	platform_green_alpha[28][29] = 1'b1; \
	platform_green_alpha[28][30] = 1'b1; \
	platform_green_alpha[28][31] = 1'b1; \
	platform_green_alpha[28][32] = 1'b1; \
	platform_green_alpha[28][33] = 1'b1; \
	platform_green_alpha[28][34] = 1'b1; \
	platform_green_alpha[28][35] = 1'b1; \
	platform_green_alpha[28][36] = 1'b1; \
	platform_green_alpha[28][37] = 1'b1; \
	platform_green_alpha[28][38] = 1'b1; \
	platform_green_alpha[28][39] = 1'b1; \
	platform_green_alpha[28][40] = 1'b1; \
	platform_green_alpha[28][41] = 1'b1; \
	platform_green_alpha[28][42] = 1'b1; \
	platform_green_alpha[28][43] = 1'b1; \
	platform_green_alpha[28][44] = 1'b1; \
	platform_green_alpha[28][45] = 1'b1; \
	platform_green_alpha[28][46] = 1'b1; \
	platform_green_alpha[28][47] = 1'b1; \
	platform_green_alpha[28][48] = 1'b1; \
	platform_green_alpha[28][49] = 1'b1; \
	platform_green_alpha[28][50] = 1'b1; \
	platform_green_alpha[28][51] = 1'b1; \
	platform_green_alpha[28][52] = 1'b1; \
	platform_green_alpha[28][53] = 1'b1; \
	platform_green_alpha[28][54] = 1'b1; \
	platform_green_alpha[28][55] = 1'b1; \
	platform_green_alpha[28][56] = 1'b1; \
	platform_green_alpha[28][57] = 1'b1; \
	platform_green_alpha[28][58] = 1'b1; \
	platform_green_alpha[28][59] = 1'b1; \
	platform_green_alpha[28][60] = 1'b1; \
	platform_green_alpha[28][61] = 1'b1; \
	platform_green_alpha[28][62] = 1'b1; \
	platform_green_alpha[28][63] = 1'b1; \
	platform_green_alpha[28][64] = 1'b1; \
	platform_green_alpha[28][65] = 1'b1; \
	platform_green_alpha[28][66] = 1'b1; \
	platform_green_alpha[28][67] = 1'b1; \
	platform_green_alpha[28][68] = 1'b1; \
	platform_green_alpha[28][69] = 1'b1; \
	platform_green_alpha[28][70] = 1'b1; \
	platform_green_alpha[28][71] = 1'b1; \
	platform_green_alpha[28][72] = 1'b1; \
	platform_green_alpha[28][73] = 1'b1; \
	platform_green_alpha[28][74] = 1'b1; \
	platform_green_alpha[28][75] = 1'b1; \
	platform_green_alpha[28][76] = 1'b1; \
	platform_green_alpha[28][77] = 1'b1; \
	platform_green_alpha[28][78] = 1'b1; \
	platform_green_alpha[28][79] = 1'b1; \
	platform_green_alpha[28][80] = 1'b1; \
	platform_green_alpha[28][81] = 1'b1; \
	platform_green_alpha[28][82] = 1'b1; \
	platform_green_alpha[28][83] = 1'b1; \
	platform_green_alpha[28][84] = 1'b1; \
	platform_green_alpha[28][85] = 1'b1; \
	platform_green_alpha[28][86] = 1'b1; \
	platform_green_alpha[28][87] = 1'b1; \
	platform_green_alpha[28][88] = 1'b1; \
	platform_green_alpha[28][89] = 1'b1; \
	platform_green_alpha[28][90] = 1'b1; \
	platform_green_alpha[28][91] = 1'b1; \
	platform_green_alpha[28][92] = 1'b1; \
	platform_green_alpha[28][93] = 1'b1; \
	platform_green_alpha[28][94] = 1'b1; \
	platform_green_alpha[28][95] = 1'b1; \
	platform_green_alpha[28][96] = 1'b1; \
	platform_green_alpha[28][97] = 1'b1; \
	platform_green_alpha[28][98] = 1'b1; \
	platform_green_alpha[28][99] = 1'b1; \
	platform_green_alpha[29][0] = 1'b1; \
	platform_green_alpha[29][1] = 1'b1; \
	platform_green_alpha[29][2] = 1'b1; \
	platform_green_alpha[29][3] = 1'b1; \
	platform_green_alpha[29][4] = 1'b1; \
	platform_green_alpha[29][5] = 1'b1; \
	platform_green_alpha[29][6] = 1'b1; \
	platform_green_alpha[29][7] = 1'b1; \
	platform_green_alpha[29][8] = 1'b1; \
	platform_green_alpha[29][9] = 1'b1; \
	platform_green_alpha[29][10] = 1'b1; \
	platform_green_alpha[29][11] = 1'b1; \
	platform_green_alpha[29][12] = 1'b1; \
	platform_green_alpha[29][13] = 1'b1; \
	platform_green_alpha[29][14] = 1'b1; \
	platform_green_alpha[29][15] = 1'b1; \
	platform_green_alpha[29][16] = 1'b1; \
	platform_green_alpha[29][17] = 1'b1; \
	platform_green_alpha[29][18] = 1'b1; \
	platform_green_alpha[29][19] = 1'b1; \
	platform_green_alpha[29][20] = 1'b1; \
	platform_green_alpha[29][21] = 1'b1; \
	platform_green_alpha[29][22] = 1'b1; \
	platform_green_alpha[29][23] = 1'b1; \
	platform_green_alpha[29][24] = 1'b1; \
	platform_green_alpha[29][25] = 1'b1; \
	platform_green_alpha[29][26] = 1'b1; \
	platform_green_alpha[29][27] = 1'b1; \
	platform_green_alpha[29][28] = 1'b1; \
	platform_green_alpha[29][29] = 1'b1; \
	platform_green_alpha[29][30] = 1'b1; \
	platform_green_alpha[29][31] = 1'b1; \
	platform_green_alpha[29][32] = 1'b1; \
	platform_green_alpha[29][33] = 1'b1; \
	platform_green_alpha[29][34] = 1'b1; \
	platform_green_alpha[29][35] = 1'b1; \
	platform_green_alpha[29][36] = 1'b1; \
	platform_green_alpha[29][37] = 1'b1; \
	platform_green_alpha[29][38] = 1'b1; \
	platform_green_alpha[29][39] = 1'b1; \
	platform_green_alpha[29][40] = 1'b1; \
	platform_green_alpha[29][41] = 1'b1; \
	platform_green_alpha[29][42] = 1'b1; \
	platform_green_alpha[29][43] = 1'b1; \
	platform_green_alpha[29][44] = 1'b1; \
	platform_green_alpha[29][45] = 1'b1; \
	platform_green_alpha[29][46] = 1'b1; \
	platform_green_alpha[29][47] = 1'b1; \
	platform_green_alpha[29][48] = 1'b1; \
	platform_green_alpha[29][49] = 1'b1; \
	platform_green_alpha[29][50] = 1'b1; \
	platform_green_alpha[29][51] = 1'b1; \
	platform_green_alpha[29][52] = 1'b1; \
	platform_green_alpha[29][53] = 1'b1; \
	platform_green_alpha[29][54] = 1'b1; \
	platform_green_alpha[29][55] = 1'b1; \
	platform_green_alpha[29][56] = 1'b1; \
	platform_green_alpha[29][57] = 1'b1; \
	platform_green_alpha[29][58] = 1'b1; \
	platform_green_alpha[29][59] = 1'b1; \
	platform_green_alpha[29][60] = 1'b1; \
	platform_green_alpha[29][61] = 1'b1; \
	platform_green_alpha[29][62] = 1'b1; \
	platform_green_alpha[29][63] = 1'b1; \
	platform_green_alpha[29][64] = 1'b1; \
	platform_green_alpha[29][65] = 1'b1; \
	platform_green_alpha[29][66] = 1'b1; \
	platform_green_alpha[29][67] = 1'b1; \
	platform_green_alpha[29][68] = 1'b1; \
	platform_green_alpha[29][69] = 1'b1; \
	platform_green_alpha[29][70] = 1'b1; \
	platform_green_alpha[29][71] = 1'b1; \
	platform_green_alpha[29][72] = 1'b1; \
	platform_green_alpha[29][73] = 1'b1; \
	platform_green_alpha[29][74] = 1'b1; \
	platform_green_alpha[29][75] = 1'b1; \
	platform_green_alpha[29][76] = 1'b1; \
	platform_green_alpha[29][77] = 1'b1; \
	platform_green_alpha[29][78] = 1'b1; \
	platform_green_alpha[29][79] = 1'b1; \
	platform_green_alpha[29][80] = 1'b1; \
	platform_green_alpha[29][81] = 1'b1; \
	platform_green_alpha[29][82] = 1'b1; \
	platform_green_alpha[29][83] = 1'b1; \
	platform_green_alpha[29][84] = 1'b1; \
	platform_green_alpha[29][85] = 1'b1; \
	platform_green_alpha[29][86] = 1'b1; \
	platform_green_alpha[29][87] = 1'b1; \
	platform_green_alpha[29][88] = 1'b1; \
	platform_green_alpha[29][89] = 1'b1; \
	platform_green_alpha[29][90] = 1'b1; \
	platform_green_alpha[29][91] = 1'b1; \
	platform_green_alpha[29][92] = 1'b1; \
	platform_green_alpha[29][93] = 1'b1; \
	platform_green_alpha[29][94] = 1'b1; \
	platform_green_alpha[29][95] = 1'b1; \
	platform_green_alpha[29][96] = 1'b1; \
	platform_green_alpha[29][97] = 1'b1; \
	platform_green_alpha[29][98] = 1'b1; \
	platform_green_alpha[29][99] = 1'b1; \
end

`endif // INITIAL_PLATFORM_GREEN
