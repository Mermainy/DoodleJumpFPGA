module platforms(
	output [4:0][3:0][1:0] platforms
);



endmodule
